module micro_ucr_hash ( gnd, vdd, clk, bloque_datos, inicio, target, bounty, terminado);

input gnd, vdd;
input clk;
input inicio;
output terminado;
input [95:0] bloque_datos;
input [7:0] target;
output [123:0] bounty;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_3917_), .Y(_3917__bF_buf4) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_3917_), .Y(_3917__bF_buf3) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_3917_), .Y(_3917__bF_buf2) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_3917_), .Y(_3917__bF_buf1) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(_3917_), .Y(_3917__bF_buf0) );
CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(_3860_), .Y(_3860__bF_buf4) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(_3860_), .Y(_3860__bF_buf3) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(_3860_), .Y(_3860__bF_buf2) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(_3860_), .Y(_3860__bF_buf1) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(_3860_), .Y(_3860__bF_buf0) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(_3777_), .Y(_3777__bF_buf4) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(_3777_), .Y(_3777__bF_buf3) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_3777_), .Y(_3777__bF_buf2) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(_3777_), .Y(_3777__bF_buf1) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(_3777_), .Y(_3777__bF_buf0) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(_3964_), .Y(_3964__bF_buf4) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(_3964_), .Y(_3964__bF_buf3) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(_3964_), .Y(_3964__bF_buf2) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(_3964_), .Y(_3964__bF_buf1) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(_3964_), .Y(_3964__bF_buf0) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_0__0_), .Y(bounty[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_0__1_), .Y(bounty[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_0__2_), .Y(bounty[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_0__3_), .Y(bounty[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(bounty[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(bounty[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(bounty[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(bounty[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(bounty[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(bounty[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(bounty[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(bounty[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(bounty[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(bounty[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(bounty[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(bounty[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(bounty[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(bounty[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(bounty[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(bounty[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(bounty[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(bounty[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(bounty[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(bounty[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[31]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[32]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[33]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[34]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[35]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[36]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[37]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[38]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[39]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[40]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[41]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[42]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[43]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[44]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[45]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[46]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[47]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[48]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[49]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[50]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[51]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[52]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[53]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[54]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[55]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[56]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[57]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[58]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[59]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[60]) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[61]) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[62]) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[63]) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[64]) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[65]) );
BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[66]) );
BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[67]) );
BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[68]) );
BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[69]) );
BUFX2 BUFX2_71 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[70]) );
BUFX2 BUFX2_72 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[71]) );
BUFX2 BUFX2_73 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[72]) );
BUFX2 BUFX2_74 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[73]) );
BUFX2 BUFX2_75 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[74]) );
BUFX2 BUFX2_76 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[75]) );
BUFX2 BUFX2_77 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[76]) );
BUFX2 BUFX2_78 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[77]) );
BUFX2 BUFX2_79 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[78]) );
BUFX2 BUFX2_80 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[79]) );
BUFX2 BUFX2_81 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[80]) );
BUFX2 BUFX2_82 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[81]) );
BUFX2 BUFX2_83 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[82]) );
BUFX2 BUFX2_84 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[83]) );
BUFX2 BUFX2_85 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[84]) );
BUFX2 BUFX2_86 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[85]) );
BUFX2 BUFX2_87 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[86]) );
BUFX2 BUFX2_88 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[87]) );
BUFX2 BUFX2_89 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[88]) );
BUFX2 BUFX2_90 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[89]) );
BUFX2 BUFX2_91 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[90]) );
BUFX2 BUFX2_92 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[91]) );
BUFX2 BUFX2_93 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[92]) );
BUFX2 BUFX2_94 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[93]) );
BUFX2 BUFX2_95 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[94]) );
BUFX2 BUFX2_96 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[95]) );
BUFX2 BUFX2_97 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[96]) );
BUFX2 BUFX2_98 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[97]) );
BUFX2 BUFX2_99 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[98]) );
BUFX2 BUFX2_100 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[99]) );
BUFX2 BUFX2_101 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[100]) );
BUFX2 BUFX2_102 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[101]) );
BUFX2 BUFX2_103 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[102]) );
BUFX2 BUFX2_104 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[103]) );
BUFX2 BUFX2_105 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[104]) );
BUFX2 BUFX2_106 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[105]) );
BUFX2 BUFX2_107 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[106]) );
BUFX2 BUFX2_108 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[107]) );
BUFX2 BUFX2_109 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[108]) );
BUFX2 BUFX2_110 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[109]) );
BUFX2 BUFX2_111 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[110]) );
BUFX2 BUFX2_112 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[111]) );
BUFX2 BUFX2_113 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[112]) );
BUFX2 BUFX2_114 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[113]) );
BUFX2 BUFX2_115 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[114]) );
BUFX2 BUFX2_116 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[115]) );
BUFX2 BUFX2_117 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[116]) );
BUFX2 BUFX2_118 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[117]) );
BUFX2 BUFX2_119 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[118]) );
BUFX2 BUFX2_120 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[119]) );
BUFX2 BUFX2_121 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[120]) );
BUFX2 BUFX2_122 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[121]) );
BUFX2 BUFX2_123 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[122]) );
BUFX2 BUFX2_124 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(bounty[123]) );
BUFX2 BUFX2_125 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(terminado) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(_503_), .Y(_867_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[22]), .B(_857_), .C(_861_), .Y(_868_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_863_), .C(_864_), .Y(_869_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_869_), .C(_867_), .Y(_870_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_866_), .B(_870_), .C(_801_), .Y(_871_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_512_), .Y(_872_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_868_), .C(_869_), .Y(_873_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_862_), .C(_865_), .Y(_874_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_873_), .C(_874_), .Y(_875_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3322_), .B(_3326_), .Y(_876_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .Y(_877_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_877_), .Y(_878_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_877_), .B(_855_), .Y(_879_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_878_), .B(_879_), .Y(_880_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_880_), .Y(_881_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_880_), .B(_320_), .Y(_882_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_882_), .B(_881_), .C(_324_), .Y(_883_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(_324_), .Y(_884_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_882_), .Y(_885_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_884_), .B(_885_), .Y(_886_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_883_), .B(_886_), .Y(_887_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_876_), .B(_887_), .Y(_888_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_888_), .B(_875_), .C(_871_), .Y(_889_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(_874_), .C(_872_), .Y(_890_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_862_), .C(_865_), .Y(_891_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_868_), .C(_869_), .Y(_892_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_892_), .C(_801_), .Y(_893_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_888_), .Y(_894_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_890_), .C(_894_), .Y(_895_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_889_), .C(_895_), .Y(_896_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_894_), .B(_875_), .C(_871_), .Y(_897_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_890_), .C(_888_), .Y(_898_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[38]), .B(_897_), .C(_898_), .Y(_899_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_896_), .B(_899_), .C(_524_), .Y(_900_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(_524_), .Y(_901_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[38]), .B(_889_), .C(_895_), .Y(_902_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_897_), .C(_898_), .Y(_903_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_902_), .B(_903_), .C(_901_), .Y(_904_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_900_), .B(_904_), .C(_799_), .Y(_905_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_533_), .Y(_906_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_902_), .C(_903_), .Y(_907_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_896_), .C(_899_), .Y(_908_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_906_), .B(_907_), .C(_908_), .Y(_909_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_3333_), .B(_3337_), .Y(_910_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[26]), .B(_883_), .C(_886_), .Y(_911_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[26]), .Y(_912_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_883_), .Y(_913_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_884_), .Y(_914_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_914_), .B(_913_), .C(_912_), .Y(_915_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_911_), .B(_915_), .C(_327_), .Y(_916_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_327_), .Y(_917_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_913_), .B(_912_), .C(_914_), .Y(_918_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_883_), .B(_886_), .C(bloque_datos[26]), .Y(_919_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_919_), .C(_918_), .Y(_920_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_920_), .B(_916_), .C(_331_), .Y(_921_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(_331_), .Y(_922_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_920_), .Y(_923_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_923_), .Y(_924_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_921_), .B(_924_), .Y(_925_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_925_), .Y(_926_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_926_), .C(_905_), .Y(_927_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_907_), .B(_908_), .C(_906_), .Y(_928_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_896_), .C(_899_), .Y(_929_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_902_), .C(_903_), .Y(_930_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_533_), .C(_929_), .D(_930_), .Y(_931_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_926_), .Y(_932_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_928_), .C(_932_), .Y(_933_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_927_), .C(_933_), .Y(_934_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_932_), .C(_905_), .Y(_935_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_928_), .C(_926_), .Y(_936_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[54]), .B(_935_), .C(_936_), .Y(_937_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_937_), .C(_545_), .Y(_938_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(_545_), .Y(_939_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[54]), .B(_927_), .C(_933_), .Y(_940_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_935_), .C(_936_), .Y(_941_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_941_), .C(_939_), .Y(_942_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_942_), .C(_797_), .Y(_943_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_554_), .Y(_944_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_939_), .B(_940_), .C(_941_), .Y(_945_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_934_), .C(_937_), .Y(_946_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(_945_), .C(_946_), .Y(_947_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_338_), .Y(_948_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[42]), .B(_921_), .C(_924_), .Y(_949_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[42]), .Y(_950_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_921_), .Y(_951_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_922_), .Y(_952_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_951_), .C(_950_), .Y(_953_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(_953_), .C(_334_), .Y(_954_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_954_), .Y(_955_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_949_), .C(_953_), .Y(_956_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_955_), .C(_948_), .Y(_957_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(_956_), .Y(_958_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_954_), .C(_958_), .Y(_959_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_957_), .B(_959_), .Y(_960_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_3349_), .B(_3346_), .C(_960_), .Y(_961_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3346_), .B(_3349_), .Y(_962_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_957_), .B(_959_), .C(_962_), .Y(_963_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_961_), .B(_963_), .Y(_964_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_964_), .C(_943_), .Y(_965_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_945_), .B(_946_), .C(_944_), .Y(_966_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_939_), .B(_934_), .C(_937_), .Y(_967_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_940_), .C(_941_), .Y(_968_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_968_), .C(_797_), .Y(_969_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_964_), .Y(_970_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(_966_), .C(_970_), .Y(_971_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_965_), .C(_971_), .Y(_972_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_966_), .B(_969_), .C(_964_), .Y(_973_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_970_), .C(_943_), .Y(_974_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[70]), .B(_974_), .C(_973_), .Y(_975_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_975_), .C(_566_), .Y(_976_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(_566_), .Y(_977_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[70]), .B(_965_), .C(_971_), .Y(_978_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_974_), .C(_973_), .Y(_979_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_979_), .C(_977_), .Y(_980_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_980_), .C(_795_), .Y(_981_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_575_), .Y(_982_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_977_), .B(_978_), .C(_979_), .Y(_983_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_972_), .C(_975_), .Y(_984_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_983_), .C(_984_), .Y(_985_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_344_), .Y(_986_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_341_), .Y(_987_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[58]), .Y(_988_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_957_), .B(_988_), .C(_959_), .Y(_989_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_958_), .B(_954_), .C(_338_), .Y(_990_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_948_), .B(_956_), .C(_955_), .Y(_991_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_991_), .C(bloque_datos[58]), .Y(_992_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_989_), .B(_992_), .C(_987_), .Y(_993_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[58]), .B(_990_), .C(_991_), .Y(_994_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_959_), .B(_957_), .C(_988_), .Y(_995_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_994_), .C(_995_), .Y(_996_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_993_), .C(_986_), .Y(_997_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_995_), .C(_341_), .Y(_998_) );
NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_987_), .B(_992_), .C(_989_), .Y(_999_) );
NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_998_), .C(_999_), .Y(_1000_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_1000_), .Y(_1001_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_3361_), .B(_3358_), .C(_1001_), .Y(_1002_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3358_), .B(_3361_), .Y(_1003_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_1000_), .C(_1003_), .Y(_1004_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1002_), .B(_1004_), .Y(_1005_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_985_), .B(_1005_), .C(_981_), .Y(_1006_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_984_), .C(_982_), .Y(_1007_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_977_), .B(_972_), .C(_975_), .Y(_1008_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_978_), .C(_979_), .Y(_1009_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_1009_), .C(_795_), .Y(_1010_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .Y(_1011_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_1007_), .C(_1011_), .Y(_1012_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_1006_), .C(_1012_), .Y(_1013_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_985_), .B(_1011_), .C(_981_), .Y(_1014_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_1007_), .C(_1005_), .Y(_1015_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[86]), .B(_1014_), .C(_1015_), .Y(_1016_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .B(_1016_), .C(_588_), .Y(_1017_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(_588_), .Y(_1018_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[86]), .B(_1006_), .C(_1012_), .Y(_1019_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_1014_), .C(_1015_), .Y(_1020_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1020_), .C(_1018_), .Y(_1021_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .B(_1021_), .C(_793_), .Y(_1022_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_597_), .Y(_1023_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1018_), .B(_1019_), .C(_1020_), .Y(_1024_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_1013_), .C(_1016_), .Y(_1025_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(_1024_), .C(_1025_), .Y(_1026_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3370_), .B(_3373_), .Y(_1027_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .Y(_1028_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_998_), .C(_344_), .Y(_1029_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_986_), .C(_993_), .Y(_1030_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[74]), .B(_1030_), .C(_1029_), .Y(_1031_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[74]), .Y(_1032_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .B(_997_), .C(_1032_), .Y(_1033_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .B(_1033_), .C(_347_), .Y(_1034_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_347_), .Y(_1035_) );
NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1032_), .B(_997_), .C(_1000_), .Y(_1036_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1030_), .B(_1029_), .C(bloque_datos[74]), .Y(_1037_) );
NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_1037_), .C(_1036_), .Y(_1038_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1038_), .B(_1034_), .C(_350_), .Y(_1039_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_349_), .Y(_1040_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1036_), .B(_1037_), .C(_1035_), .Y(_1041_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_1031_), .C(_1033_), .Y(_1042_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1042_), .B(_1040_), .C(_1041_), .Y(_1043_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1043_), .C(_1028_), .Y(_1044_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1043_), .B(_1039_), .Y(_1045_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(_1027_), .Y(_1046_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_1044_), .Y(_1047_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .B(_1047_), .C(_1022_), .Y(_1048_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1024_), .B(_1025_), .C(_1023_), .Y(_1049_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1018_), .B(_1013_), .C(_1016_), .Y(_1050_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_1019_), .C(_1020_), .Y(_1051_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1050_), .B(_1051_), .C(_793_), .Y(_1052_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_1047_), .Y(_1053_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1052_), .B(_1049_), .C(_1053_), .Y(_1054_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_1048_), .C(_1054_), .Y(_1055_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .B(_1053_), .C(_1022_), .Y(_1056_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1052_), .B(_1049_), .C(_1047_), .Y(_1057_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(W_134_), .B(_1056_), .C(_1057_), .Y(_1058_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1058_), .C(_609_), .Y(_1059_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(_609_), .Y(_1060_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(W_134_), .B(_1048_), .C(_1054_), .Y(_1061_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_1056_), .C(_1057_), .Y(_1062_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_1062_), .C(_1060_), .Y(_1063_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .B(_1063_), .C(_791_), .Y(_1064_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_618_), .Y(_1065_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1060_), .B(_1061_), .C(_1062_), .Y(_1066_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_1055_), .C(_1058_), .Y(_1067_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1065_), .B(_1066_), .C(_1067_), .Y(_1068_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(bloque_datos[90]), .Y(_1069_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_1069_), .Y(_1070_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .B(_354_), .Y(_1071_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1071_), .B(_1070_), .C(_358_), .Y(_1072_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .B(_1071_), .Y(_1073_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_1073_), .Y(_1074_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_1074_), .Y(_1075_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1075_), .C(_1064_), .Y(_1076_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_1067_), .C(_1065_), .Y(_1077_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1060_), .B(_1055_), .C(_1058_), .Y(_1078_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_1061_), .C(_1062_), .Y(_1079_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1078_), .B(_1079_), .C(_791_), .Y(_1080_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_1074_), .B(_1072_), .Y(_1081_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1077_), .C(_1081_), .Y(_1082_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_1076_), .C(_1082_), .Y(_1083_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_1083_), .Y(_1084_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1077_), .C(_1075_), .Y(_1085_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1081_), .C(_1064_), .Y(_1086_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1086_), .B(_1085_), .C(_789_), .Y(_1087_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(W_150_), .B(_1087_), .Y(_1088_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_1084_), .C(_1088_), .Y(_1089_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(W_150_), .B(_1083_), .Y(_1090_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_1087_), .Y(_1091_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_1090_), .C(_1091_), .Y(_1092_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_1089_), .C(_1092_), .Y(_1093_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_640_), .Y(_1094_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_1090_), .C(_1091_), .Y(_1095_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_1084_), .C(_1088_), .Y(_1096_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1094_), .B(_1096_), .C(_1095_), .Y(_1097_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(W_138_), .B(_1081_), .Y(_1098_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(W_138_), .Y(_1099_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1099_), .B(_1075_), .Y(_1100_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1100_), .B(_1098_), .Y(_1101_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .B(_362_), .Y(_1102_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_365_), .C(_1102_), .Y(_1103_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_367_), .Y(_1104_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1103_), .B(_1104_), .Y(_1105_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(_1093_), .C(_1097_), .Y(_1106_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .B(_1095_), .C(_1094_), .Y(_1107_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_1092_), .C(_787_), .Y(_1108_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .Y(_1109_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1107_), .B(_1108_), .C(_1109_), .Y(_1110_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_1106_), .C(_1110_), .Y(_1111_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_1111_), .Y(_1112_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1107_), .B(_1108_), .C(_1105_), .Y(_1113_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1109_), .B(_1093_), .C(_1097_), .Y(_1114_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1114_), .B(_1113_), .C(_784_), .Y(_1115_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(W_166_), .B(_1115_), .Y(_1116_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_1112_), .C(_1116_), .Y(_1117_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(W_166_), .B(_1111_), .Y(_1118_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_1115_), .Y(_1119_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_651_), .B(_1118_), .C(_1119_), .Y(_1120_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(_1117_), .C(_1120_), .Y(_1121_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_656_), .Y(_1122_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_1118_), .C(_1119_), .Y(_1123_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_651_), .B(_1112_), .C(_1116_), .Y(_1124_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_1124_), .C(_1122_), .Y(_1125_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(W_154_), .Y(_1126_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1126_), .B(_1105_), .Y(_1127_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(W_154_), .B(_1109_), .Y(_1128_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(_1127_), .C(_371_), .Y(_1129_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_1129_), .Y(_1130_) );
NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_1127_), .C(_1128_), .Y(_1131_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1131_), .C(_374_), .Y(_1132_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_374_), .Y(_1133_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_1131_), .Y(_1134_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .B(_1129_), .C(_1134_), .Y(_1135_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .B(_1135_), .Y(_1136_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1136_), .C(_1125_), .Y(_1137_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_1124_), .C(_1122_), .Y(_1138_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1117_), .B(_1120_), .C(_782_), .Y(_1139_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_1132_), .Y(_1140_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(_1139_), .C(_1140_), .Y(_1141_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_1137_), .C(_1141_), .Y(_1142_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_1142_), .Y(_1143_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1140_), .C(_1125_), .Y(_1144_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(_1139_), .C(_1136_), .Y(_1145_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .B(_1145_), .Y(_1146_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(W_182_), .B(_780_), .C(_1146_), .Y(_1147_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_1147_), .C(_1143_), .Y(_1148_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(W_182_), .B(_1142_), .Y(_1149_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_780_), .C(_1146_), .Y(_1150_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_1150_), .C(_1149_), .Y(_1151_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_1148_), .C(_1151_), .Y(_1152_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_674_), .Y(_1153_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_676_), .C(_671_), .Y(_1154_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_1150_), .C(_1149_), .Y(_1155_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_1147_), .C(_1143_), .Y(_1156_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_1156_), .C(_1154_), .Y(_1157_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_379_), .Y(_1158_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(W_170_), .Y(_1159_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(W_170_), .B(_1140_), .Y(_1160_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(_1160_), .C(_1158_), .Y(_1161_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_1161_), .Y(_1162_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_1159_), .Y(_1163_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_379_), .Y(_1164_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1164_), .B(_1162_), .C(_383_), .Y(_1165_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_383_), .Y(_1166_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_1163_), .Y(_1167_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1166_), .B(_1161_), .C(_1167_), .Y(_1168_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1168_), .B(_1165_), .Y(_1169_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1152_), .C(_1157_), .Y(_1170_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_1156_), .C(_1154_), .Y(_1171_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1148_), .B(_1151_), .C(_777_), .Y(_1172_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(_1168_), .Y(_1173_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1171_), .B(_1172_), .C(_1173_), .Y(_1174_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_775_), .B(_1170_), .C(_1174_), .Y(_1175_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_1175_), .Y(_1176_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1171_), .B(_1172_), .C(_1169_), .Y(_1177_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1173_), .B(_1152_), .C(_1157_), .Y(_1178_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(_1177_), .Y(_1179_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(W_198_), .B(_775_), .C(_1179_), .Y(_1180_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(_1176_), .C(_1180_), .Y(_1181_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(W_198_), .B(_1175_), .Y(_1182_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(_1177_), .C(_774_), .Y(_1183_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_1183_), .Y(_1184_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_1182_), .C(_1184_), .Y(_1185_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_1181_), .C(_1185_), .Y(_1186_) );
NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_427_), .C(_689_), .Y(_1187_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(_695_), .C(_690_), .Y(_1188_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(_1182_), .C(_1184_), .Y(_1189_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_1176_), .C(_1180_), .Y(_1190_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1188_), .B(_1190_), .C(_1189_), .Y(_1191_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(_391_), .Y(_1192_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_387_), .Y(_1193_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(W_186_), .Y(_1194_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1194_), .B(_1169_), .Y(_1195_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(W_186_), .B(_1173_), .Y(_1196_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1196_), .B(_1195_), .C(_1193_), .Y(_1197_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1196_), .Y(_1198_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_1198_), .Y(_1199_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(_1199_), .Y(_1200_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1200_), .B(_1192_), .Y(_1201_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .Y(_1202_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_1191_), .C(_1202_), .Y(_1203_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1202_), .B(_1186_), .C(_1191_), .Y(_1204_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_3428_), .B(_3432_), .C(_1204_), .Y(_1205_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(_1203_), .C(_770_), .Y(_1206_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_1191_), .Y(_1207_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .B(_1207_), .Y(_1208_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(_3437_), .Y(_1209_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_1204_), .B(_1209_), .Y(_1210_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(W_214_), .B(_1208_), .C(_1210_), .Y(_1211_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1206_), .B(_1211_), .C(_708_), .Y(_1212_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(_1203_), .C(W_214_), .Y(_1213_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_770_), .B(_1208_), .C(_1210_), .Y(_1214_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1213_), .B(_1214_), .C(_711_), .Y(_1215_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1212_), .B(_1215_), .C(_769_), .Y(_1216_) );
NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_424_), .C(_708_), .Y(_1217_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1217_), .B(_714_), .C(_709_), .Y(_1218_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_1213_), .C(_1214_), .Y(_1219_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_1206_), .C(_1211_), .Y(_1220_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1219_), .B(_1220_), .C(_1218_), .Y(_1221_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(_395_), .Y(_1222_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(W_202_), .B(_1201_), .Y(_1223_) );
INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .Y(_1224_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(W_202_), .B(_1201_), .Y(_1225_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .B(_1225_), .C(_1222_), .Y(_1226_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .Y(_1227_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .B(_1225_), .Y(_1228_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .B(_1228_), .Y(_1229_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1229_), .B(_1227_), .C(_399_), .Y(_1230_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_399_), .Y(_1231_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_1222_), .Y(_1232_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1231_), .B(_1226_), .C(_1232_), .Y(_1233_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1230_), .B(_1233_), .Y(_1234_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .B(_1234_), .C(_1216_), .Y(_1235_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1219_), .B(_1220_), .C(_1218_), .Y(_1236_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_1206_), .C(_1211_), .Y(_1237_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_1213_), .C(_1214_), .Y(_1238_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1238_), .B(_1237_), .C(_769_), .Y(_1239_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_1233_), .B(_1230_), .Y(_1240_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_1239_), .C(_1240_), .Y(_1241_) );
NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_1235_), .C(_1241_), .Y(_1242_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_765_), .B(_1242_), .Y(_1243_) );
NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .B(_1240_), .C(_1216_), .Y(_1244_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_1239_), .C(_1234_), .Y(_1245_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .B(_1245_), .C(_766_), .Y(_1246_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(W_230_), .B(_1246_), .Y(_1247_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1243_), .B(_1247_), .C(_727_), .Y(_1248_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(W_230_), .B(_1242_), .Y(_1249_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_765_), .B(_1246_), .Y(_1250_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1249_), .B(_1250_), .C(_730_), .Y(_1251_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1248_), .B(_1251_), .C(_764_), .Y(_1252_) );
NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_723_), .B(_421_), .C(_727_), .Y(_1253_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1253_), .B(_733_), .C(_728_), .Y(_1254_) );
NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_730_), .B(_1249_), .C(_1250_), .Y(_1255_) );
NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_1243_), .C(_1247_), .Y(_1256_) );
NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_1255_), .C(_1254_), .Y(_1257_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(W_218_), .B(_1240_), .Y(_1258_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(W_218_), .Y(_1259_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1259_), .B(_1234_), .Y(_1260_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1260_), .B(_1258_), .C(_403_), .Y(_1261_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_403_), .Y(_1262_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1260_), .B(_1258_), .Y(_1263_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1262_), .B(_1263_), .Y(_1264_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .B(_1261_), .C(_407_), .Y(_1265_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_407_), .Y(_1266_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .Y(_1267_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_1263_), .B(_1262_), .Y(_1268_) );
NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_1267_), .C(_1268_), .Y(_1269_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .B(_1269_), .Y(_1270_) );
NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1270_), .B(_1257_), .C(_1252_), .Y(_1271_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_1255_), .C(_1254_), .Y(_1272_) );
NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_730_), .B(_1243_), .C(_1247_), .Y(_1273_) );
NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_1249_), .C(_1250_), .Y(_1274_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1273_), .B(_1274_), .C(_764_), .Y(_1275_) );
INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(_1270_), .Y(_1276_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .B(_1275_), .C(_1276_), .Y(_1277_) );
NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_3457_), .B(_1271_), .C(_1277_), .Y(_1278_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(W_246_), .B(_1278_), .Y(_1279_) );
INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(W_246_), .Y(_1280_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .B(_1275_), .C(_1270_), .Y(_1281_) );
NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_1257_), .C(_1252_), .Y(_1282_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1282_), .B(_1281_), .C(_3456_), .Y(_1283_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_1283_), .Y(_1284_) );
NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(_744_), .B(_1279_), .C(_1284_), .Y(_1285_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_1278_), .Y(_1286_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(W_246_), .B(_1283_), .Y(_1287_) );
NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_748_), .B(_1286_), .C(_1287_), .Y(_1288_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1285_), .B(_1288_), .C(_762_), .Y(_1289_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_753_), .C(_745_), .Y(_1290_) );
NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_744_), .B(_1286_), .C(_1287_), .Y(_1291_) );
NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_748_), .B(_1279_), .C(_1284_), .Y(_1292_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1291_), .B(_1292_), .C(_1290_), .Y(_1293_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(W_234_), .B(_1276_), .Y(_1294_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(W_234_), .Y(_1295_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1270_), .Y(_1296_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1296_), .B(_1294_), .C(_411_), .Y(_1297_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_411_), .Y(_1298_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1296_), .B(_1294_), .Y(_1299_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1298_), .B(_1299_), .Y(_1300_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1300_), .B(_1297_), .C(_415_), .Y(_1301_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_415_), .Y(_1302_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_1297_), .Y(_1303_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_1298_), .Y(_1304_) );
NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1302_), .B(_1303_), .C(_1304_), .Y(_1305_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1301_), .B(_1305_), .Y(_1306_) );
INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .Y(_1307_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1293_), .C(_1307_), .Y(_1308_) );
NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .B(_1291_), .C(_1292_), .Y(_1309_) );
NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1285_), .B(_1288_), .C(_762_), .Y(_1310_) );
NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(_1306_), .C(_1310_), .Y(_1311_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1311_), .B(_1308_), .Y(_1312_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(_759_), .Y(H_6_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1293_), .C(_1306_), .Y(_1313_) );
NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(_1307_), .C(_1310_), .Y(_1314_) );
NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(_1313_), .C(_759_), .Y(_1315_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1279_), .B(_1284_), .C(_744_), .Y(_1316_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(_1290_), .C(_1285_), .Y(_1317_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1297_), .B(_415_), .C(_1304_), .Y(_1318_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_1267_), .C(_1264_), .Y(_1319_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .Y(_1320_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1231_), .B(_1226_), .C(_1229_), .Y(_1321_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1200_), .B(_391_), .C(_1199_), .Y(_1322_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1166_), .B(_1161_), .C(_1164_), .Y(_1323_) );
INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .Y(_1324_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(W_171_), .Y(_1325_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .B(_1129_), .C(_1131_), .Y(_1326_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_360_), .C(_1101_), .Y(_1327_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_1101_), .Y(_1328_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_1327_), .C(_1328_), .Y(_1329_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_1098_), .Y(_1330_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_1073_), .C(_1071_), .Y(_1331_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[90]), .Y(_1332_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1332_), .B(_1045_), .Y(_1333_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_1034_), .C(_1042_), .Y(_1334_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[75]), .Y(_1335_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_344_), .C(_996_), .Y(_1336_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[59]), .Y(_1337_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_954_), .B(_338_), .C(_956_), .Y(_1338_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[43]), .Y(_1339_) );
NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_911_), .C(_915_), .Y(_1340_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_331_), .C(_1340_), .Y(_1341_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[27]), .Y(_1342_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_880_), .Y(_1343_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_324_), .C(_1343_), .Y(_1344_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_878_), .Y(_1345_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .Y(_1346_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_851_), .Y(_1347_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_317_), .C(_1347_), .Y(_1348_) );
INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(_848_), .Y(_1349_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(W_27_), .B(W_11_), .Y(_1350_) );
INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .Y(_1351_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(W_27_), .B(W_11_), .Y(_1352_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .B(_1351_), .Y(_1353_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1353_), .B(_1349_), .Y(_1354_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_1354_), .Y(_1355_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1346_), .B(_1355_), .Y(_1356_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1349_), .B(_1353_), .Y(_1357_) );
AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .B(_1351_), .C(_848_), .Y(_1358_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(_1357_), .Y(_1359_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_1359_), .Y(_1360_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .B(_1360_), .Y(_1361_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1361_), .B(_1356_), .Y(_1362_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_1362_), .B(_1345_), .Y(_1363_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1345_), .B(_1362_), .Y(_1364_) );
NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_1364_), .C(_1344_), .Y(_1365_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_879_), .B(_878_), .Y(_1366_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_319_), .C(_1366_), .Y(_1367_) );
AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1367_), .B(_884_), .C(_882_), .Y(_1368_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .Y(_1369_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_1364_), .Y(_1370_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1369_), .B(_1370_), .C(_1368_), .Y(_1371_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1365_), .B(_1371_), .Y(_1372_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1342_), .B(_1372_), .Y(_1373_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_1371_), .B(_1365_), .Y(_1374_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[27]), .B(_1374_), .Y(_1375_) );
NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_911_), .B(_1373_), .C(_1375_), .Y(_1376_) );
AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .B(_1375_), .C(_911_), .Y(_1377_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_1377_), .Y(_1378_) );
NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1376_), .B(_1378_), .C(_1341_), .Y(_1379_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_918_), .B(_919_), .C(_917_), .Y(_1380_) );
AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_1380_), .C(_920_), .Y(_1381_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1342_), .B(_1374_), .Y(_1382_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[27]), .B(_1372_), .Y(_1383_) );
AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1383_), .B(_1382_), .C(_918_), .Y(_1384_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1384_), .B(_1377_), .C(_1381_), .Y(_1385_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1385_), .B(_1379_), .Y(_1386_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1339_), .B(_1386_), .Y(_1387_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_1379_), .B(_1385_), .Y(_1388_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[43]), .B(_1388_), .Y(_1389_) );
NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(_1387_), .C(_1389_), .Y(_1390_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_1390_), .Y(_1391_) );
AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1387_), .B(_1389_), .C(_949_), .Y(_1392_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1392_), .B(_1391_), .Y(_1393_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_1393_), .B(_1338_), .Y(_1394_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .Y(_1395_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1391_), .B(_1392_), .C(_1395_), .Y(_1396_) );
INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(_1396_), .Y(_1397_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1394_), .B(_1397_), .C(_1337_), .Y(_1398_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_958_), .B(_959_), .C(_1393_), .Y(_1399_) );
NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[59]), .B(_1396_), .C(_1399_), .Y(_1400_) );
NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_1400_), .C(_1398_), .Y(_1401_) );
NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1337_), .B(_1396_), .C(_1399_), .Y(_1402_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1394_), .B(_1397_), .C(bloque_datos[59]), .Y(_1403_) );
NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_989_), .B(_1402_), .C(_1403_), .Y(_1404_) );
NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1401_), .C(_1404_), .Y(_1405_) );
AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1401_), .B(_1404_), .C(_1336_), .Y(_1406_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_1406_), .Y(_1407_) );
NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1335_), .B(_1405_), .C(_1407_), .Y(_1408_) );
INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(_1405_), .Y(_1409_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1409_), .B(_1406_), .C(bloque_datos[75]), .Y(_1410_) );
AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .B(_1410_), .C(_1036_), .Y(_1411_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_1411_), .Y(_1412_) );
NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1036_), .B(_1408_), .C(_1410_), .Y(_1413_) );
NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1334_), .B(_1413_), .C(_1412_), .Y(_1414_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_1334_), .Y(_1415_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_1413_), .Y(_1416_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .B(_1411_), .C(_1415_), .Y(_1417_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(_1417_), .Y(_1418_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(bloque_datos[91]), .Y(_1419_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .Y(_1420_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .Y(_1421_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1421_), .B(_1420_), .C(bloque_datos[91]), .Y(_1422_) );
AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(_1419_), .C(_1333_), .Y(_1423_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .Y(_1424_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[91]), .Y(_1425_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1421_), .B(_1420_), .C(_1425_), .Y(_1426_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(_1425_), .Y(_1427_) );
AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(_1427_), .C(_1424_), .Y(_1428_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1423_), .B(_1428_), .C(_1331_), .Y(_1429_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_1071_), .Y(_1430_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_1070_), .C(_1430_), .Y(_1431_) );
NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1424_), .B(_1426_), .C(_1427_), .Y(_1432_) );
NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .B(_1422_), .C(_1419_), .Y(_1433_) );
NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1432_), .B(_1433_), .C(_1431_), .Y(_1434_) );
NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(W_139_), .B(_1434_), .C(_1429_), .Y(_1435_) );
AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_1429_), .C(W_139_), .Y(_1436_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .Y(_1437_) );
AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1435_), .B(_1437_), .C(_1330_), .Y(_1438_) );
INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(_1435_), .Y(_1439_) );
NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1098_), .B(_1436_), .C(_1439_), .Y(_1440_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1438_), .B(_1440_), .C(_1329_), .Y(_1441_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_1441_), .Y(_1442_) );
NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1438_), .B(_1440_), .C(_1329_), .Y(_1443_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1443_), .B(_1442_), .Y(_1444_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(W_155_), .B(_1444_), .Y(_1445_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(W_155_), .Y(_1446_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1442_), .B(_1443_), .C(_1446_), .Y(_1447_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .B(_1445_), .Y(_1448_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1126_), .B(_1105_), .C(_1448_), .Y(_1449_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_1449_), .Y(_1450_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_1448_), .Y(_1451_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_1451_), .B(_1127_), .Y(_1452_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1452_), .B(_1450_), .C(_1326_), .Y(_1453_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_1326_), .Y(_1454_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_1452_), .Y(_1455_) );
NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1449_), .B(_1455_), .C(_1454_), .Y(_1456_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1453_), .B(_1456_), .Y(_1457_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1325_), .B(_1457_), .Y(_1458_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1325_), .B(_1457_), .Y(_1459_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_1459_), .Y(_1460_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1460_), .B(_1458_), .C(_1324_), .Y(_1461_) );
INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(_1461_), .Y(_1462_) );
INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(_1457_), .Y(_1463_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(W_171_), .B(_1463_), .Y(_1464_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1459_), .B(_1464_), .Y(_1465_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1324_), .B(_1465_), .Y(_1466_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_1462_), .C(_1323_), .Y(_1467_) );
INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(_1467_), .Y(_1468_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1162_), .B(_383_), .C(_1167_), .Y(_1469_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1462_), .B(_1466_), .Y(_1470_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_1470_), .B(_1469_), .Y(_1471_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(_1471_), .Y(_1472_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(W_187_), .B(_1472_), .Y(_1473_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(W_187_), .Y(_1474_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .B(_1468_), .C(_1474_), .Y(_1475_) );
AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1475_), .B(_1473_), .C(_1195_), .Y(_1476_) );
INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(_1476_), .Y(_1477_) );
NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1475_), .C(_1473_), .Y(_1478_) );
AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1477_), .B(_1478_), .C(_1322_), .Y(_1479_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_1199_), .Y(_1480_) );
AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1192_), .B(_1197_), .C(_1480_), .Y(_1481_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1478_), .B(_1477_), .Y(_1482_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1481_), .B(_1482_), .Y(_1483_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1479_), .B(_1483_), .Y(_1484_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(W_203_), .B(_1484_), .Y(_1485_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(W_203_), .Y(_1486_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1483_), .B(_1479_), .C(_1486_), .Y(_1487_) );
AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1487_), .B(_1485_), .C(_1224_), .Y(_1488_) );
NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .B(_1487_), .C(_1485_), .Y(_1489_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_1489_), .Y(_1490_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1490_), .B(_1488_), .C(_1321_), .Y(_1491_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_1488_), .Y(_1492_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1489_), .B(_1492_), .Y(_1493_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_1321_), .Y(_1494_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1491_), .B(_1494_), .Y(_1495_) );
INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(_1495_), .Y(_1496_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(W_219_), .B(_1496_), .Y(_1497_) );
AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1491_), .B(_1494_), .C(W_219_), .Y(_1498_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_1498_), .Y(_1499_) );
AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1499_), .B(_1497_), .C(_1320_), .Y(_1500_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(W_219_), .Y(_1501_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1501_), .B(_1495_), .Y(_1502_) );
NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1498_), .B(_1258_), .C(_1502_), .Y(_1503_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1500_), .B(_1503_), .C(_1319_), .Y(_1504_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .B(_407_), .C(_1268_), .Y(_1505_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_1498_), .C(_1258_), .Y(_1506_) );
NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(_1499_), .C(_1497_), .Y(_1507_) );
NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .B(_1506_), .C(_1507_), .Y(_1508_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1508_), .B(_1504_), .Y(_1509_) );
INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .Y(_1510_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(W_235_), .B(_1510_), .Y(_1511_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(W_235_), .Y(_1512_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1512_), .B(_1509_), .Y(_1513_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(W_234_), .B(_1276_), .C(_1511_), .D(_1513_), .Y(_1514_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_1514_), .Y(_1515_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1513_), .B(_1511_), .Y(_1516_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_1516_), .B(_1294_), .Y(_1517_) );
NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1318_), .B(_1515_), .C(_1517_), .Y(_1518_) );
AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1302_), .B(_1303_), .C(_1300_), .Y(_1519_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .B(_1516_), .Y(_1520_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1520_), .B(_1514_), .C(_1519_), .Y(_1521_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(_1518_), .Y(_1522_) );
AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .B(_1218_), .C(_1212_), .Y(_1523_) );
AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1182_), .B(_1184_), .C(_692_), .Y(_1524_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_772_), .C(_1189_), .Y(_1525_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .Y(_1526_) );
AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1154_), .B(_1156_), .C(_1526_), .Y(_1527_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .B(_1468_), .Y(_1528_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .Y(_1529_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .Y(_1530_) );
AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1094_), .B(_1096_), .C(_1530_), .Y(_1531_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_1444_), .Y(_1532_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .Y(_1533_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_1429_), .Y(_1534_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .Y(_1535_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1535_), .B(_1534_), .Y(_1536_) );
AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(_1025_), .C(_1017_), .Y(_1537_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_1537_), .Y(_1538_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .Y(_1539_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_795_), .B(_980_), .C(_983_), .Y(_1540_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1406_), .B(_1409_), .Y(_1541_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .Y(_1542_) );
AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(_946_), .C(_938_), .Y(_1543_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1397_), .B(_1394_), .Y(_1544_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .Y(_1545_) );
AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_906_), .B(_908_), .C(_900_), .Y(_1546_) );
AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_874_), .C(_866_), .Y(_1547_) );
AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_842_), .C(_834_), .Y(_1548_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_806_), .C(_816_), .Y(_1549_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(W_22_), .B(_813_), .Y(_1550_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_3503_), .B(_3507_), .Y(_1551_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(W_7_), .B(W_23_), .Y(_1552_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1551_), .B(_1552_), .Y(_1553_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(W_5_), .C(W_6_), .Y(_1554_) );
XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1554_), .B(W_11_), .Y(_1555_) );
XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1555_), .Y(_1556_) );
XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1550_), .B(_1556_), .Y(_1557_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_1557_), .Y(_1558_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_3516_), .B(_3514_), .Y(_1559_) );
XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1559_), .B(bloque_datos[7]), .Y(_1560_) );
XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1560_), .B(_1558_), .Y(_1561_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1549_), .B(_1561_), .Y(_1562_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(_1549_), .Y(_1563_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[23]), .Y(_1564_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_3525_), .B(_3529_), .C(_1564_), .Y(_1565_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_3529_), .B(_3525_), .Y(_1566_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[23]), .B(_1566_), .Y(_1567_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1565_), .B(_1567_), .Y(_1568_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .B(_1563_), .C(_1568_), .Y(_1569_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(_1549_), .Y(_1570_) );
NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1565_), .B(_1567_), .C(_1570_), .Y(_1571_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .B(_1569_), .Y(_1572_) );
XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_836_), .B(_1355_), .Y(_1573_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1573_), .B(_1572_), .Y(_1574_) );
XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_836_), .B(_1360_), .Y(_1575_) );
AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .B(_1571_), .C(_1575_), .Y(_1576_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1574_), .B(_1576_), .C(_1548_), .Y(_1577_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .Y(_1578_) );
NAND3X1 NAND3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .B(_1571_), .C(_1575_), .Y(_1579_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1573_), .B(_1572_), .Y(_1580_) );
NAND3X1 NAND3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1579_), .B(_1580_), .C(_1578_), .Y(_1581_) );
NAND3X1 NAND3X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .B(_1581_), .C(_1577_), .Y(_1582_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1574_), .B(_1576_), .C(_1578_), .Y(_1583_) );
NAND3X1 NAND3X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(_1579_), .C(_1580_), .Y(_1584_) );
NAND3X1 NAND3X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .B(_1584_), .C(_1583_), .Y(_1585_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .B(_1585_), .Y(_1586_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_3543_), .B(_3540_), .Y(_1587_) );
XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .B(bloque_datos[39]), .Y(_1588_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_1588_), .Y(_1589_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_1588_), .B(_868_), .Y(_1590_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1590_), .B(_1589_), .C(_1586_), .Y(_1591_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .B(_1585_), .Y(_1592_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_1588_), .B(_868_), .Y(_1593_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_1588_), .Y(_1594_) );
NAND3X1 NAND3X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1593_), .B(_1594_), .C(_1592_), .Y(_1595_) );
NAND3X1 NAND3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1547_), .B(_1591_), .C(_1595_), .Y(_1596_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_801_), .B(_870_), .C(_873_), .Y(_1597_) );
AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1593_), .B(_1594_), .C(_1592_), .Y(_1598_) );
NOR3X1 NOR3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1590_), .B(_1589_), .C(_1586_), .Y(_1599_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1598_), .B(_1599_), .C(_1597_), .Y(_1600_) );
NAND3X1 NAND3X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1386_), .B(_1596_), .C(_1600_), .Y(_1601_) );
NAND3X1 NAND3X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1597_), .B(_1591_), .C(_1595_), .Y(_1602_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1598_), .B(_1599_), .C(_1547_), .Y(_1603_) );
NAND3X1 NAND3X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1388_), .B(_1602_), .C(_1603_), .Y(_1604_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_1601_), .B(_1604_), .Y(_1605_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .B(_3557_), .C(bloque_datos[55]), .Y(_1606_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[55]), .Y(_1607_) );
NAND3X1 NAND3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1607_), .B(_3556_), .C(_3552_), .Y(_1608_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .B(_1606_), .Y(_1609_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_902_), .B(_1609_), .Y(_1610_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .B(_902_), .Y(_1611_) );
AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1610_), .B(_1611_), .C(_1605_), .Y(_1612_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1601_), .B(_1604_), .Y(_1613_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .B(_902_), .Y(_1614_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_902_), .B(_1609_), .Y(_1615_) );
NOR3X1 NOR3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1614_), .C(_1613_), .Y(_1616_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1612_), .B(_1616_), .C(_1546_), .Y(_1617_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_799_), .B(_904_), .C(_907_), .Y(_1618_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1614_), .C(_1613_), .Y(_1619_) );
NAND3X1 NAND3X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1610_), .B(_1611_), .C(_1605_), .Y(_1620_) );
NAND3X1 NAND3X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1618_), .B(_1619_), .C(_1620_), .Y(_1621_) );
NAND3X1 NAND3X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1545_), .B(_1621_), .C(_1617_), .Y(_1622_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1612_), .B(_1616_), .C(_1618_), .Y(_1623_) );
NAND3X1 NAND3X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1546_), .B(_1619_), .C(_1620_), .Y(_1624_) );
NAND3X1 NAND3X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .B(_1624_), .C(_1623_), .Y(_1625_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_1622_), .B(_1625_), .Y(_1626_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_3565_), .B(_3571_), .Y(_1627_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .B(bloque_datos[71]), .Y(_1628_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_1628_), .Y(_1629_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1628_), .B(_940_), .Y(_1630_) );
AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1630_), .B(_1629_), .C(_1626_), .Y(_1631_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .B(_1622_), .Y(_1632_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1628_), .B(_940_), .Y(_1633_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_1628_), .Y(_1634_) );
NOR3X1 NOR3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1633_), .C(_1632_), .Y(_1635_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(_1631_), .C(_1543_), .Y(_1636_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(_942_), .C(_945_), .Y(_1637_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1633_), .C(_1632_), .Y(_1638_) );
NAND3X1 NAND3X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(_1630_), .C(_1626_), .Y(_1639_) );
NAND3X1 NAND3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .B(_1638_), .C(_1639_), .Y(_1640_) );
NAND3X1 NAND3X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1542_), .B(_1640_), .C(_1636_), .Y(_1641_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(_1631_), .C(_1637_), .Y(_1642_) );
NAND3X1 NAND3X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1543_), .B(_1638_), .C(_1639_), .Y(_1643_) );
NAND3X1 NAND3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(_1643_), .C(_1642_), .Y(_1644_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .B(_1644_), .Y(_1645_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(_3581_), .Y(_1646_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1646_), .B(bloque_datos[87]), .Y(_1647_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_1647_), .Y(_1648_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(_978_), .Y(_1649_) );
NAND3X1 NAND3X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .B(_1645_), .C(_1648_), .Y(_1650_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .B(_1644_), .Y(_1651_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(_978_), .Y(_1652_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_1647_), .Y(_1653_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_1652_), .C(_1651_), .Y(_1654_) );
NAND3X1 NAND3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1650_), .B(_1540_), .C(_1654_), .Y(_1655_) );
AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_984_), .C(_976_), .Y(_1656_) );
NOR3X1 NOR3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_1652_), .C(_1651_), .Y(_1657_) );
AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .B(_1648_), .C(_1645_), .Y(_1658_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .B(_1658_), .C(_1656_), .Y(_1659_) );
AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1659_), .C(_1539_), .Y(_1660_) );
NAND3X1 NAND3X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1656_), .B(_1650_), .C(_1654_), .Y(_1661_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .B(_1658_), .C(_1540_), .Y(_1662_) );
AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1661_), .B(_1662_), .C(_1418_), .Y(_1663_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1663_), .Y(_1664_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_3588_), .B(_3591_), .Y(_1665_) );
XNOR2X1 XNOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .B(W_135_), .Y(_1666_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1666_), .Y(_1667_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1666_), .B(_1019_), .Y(_1668_) );
NAND3X1 NAND3X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1668_), .B(_1667_), .C(_1664_), .Y(_1669_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1663_), .Y(_1670_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1666_), .B(_1019_), .Y(_1671_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1666_), .Y(_1672_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1672_), .B(_1671_), .C(_1670_), .Y(_1673_) );
NAND3X1 NAND3X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1669_), .B(_1673_), .C(_1538_), .Y(_1674_) );
NOR3X1 NOR3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1671_), .B(_1672_), .C(_1670_), .Y(_1675_) );
AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1668_), .B(_1667_), .C(_1664_), .Y(_1676_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1675_), .B(_1676_), .C(_1537_), .Y(_1677_) );
AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1674_), .B(_1677_), .C(_1536_), .Y(_1678_) );
INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(_1536_), .Y(_1679_) );
NAND3X1 NAND3X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1537_), .B(_1673_), .C(_1669_), .Y(_1680_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1675_), .B(_1676_), .C(_1538_), .Y(_1681_) );
AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1680_), .B(_1681_), .C(_1679_), .Y(_1682_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1678_), .B(_1682_), .C(_1533_), .Y(_1683_) );
NAND3X1 NAND3X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1679_), .B(_1680_), .C(_1681_), .Y(_1684_) );
NAND3X1 NAND3X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1536_), .B(_1674_), .C(_1677_), .Y(_1685_) );
NAND3X1 NAND3X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_1684_), .C(_1685_), .Y(_1686_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_1683_), .B(_1686_), .Y(_1687_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .B(_1080_), .C(_1687_), .Y(_1688_) );
AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1065_), .B(_1067_), .C(_1059_), .Y(_1689_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1686_), .B(_1683_), .Y(_1690_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_3598_), .B(_3602_), .C(_1690_), .D(_1689_), .Y(_1691_) );
NAND3X1 NAND3X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_1691_), .C(_1688_), .Y(_1692_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1689_), .B(_1690_), .Y(_1693_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_791_), .B(_1063_), .C(_1066_), .Y(_1694_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1687_), .B(_1694_), .C(_3603_), .Y(_1695_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1695_), .B(_1693_), .C(_1444_), .Y(_1696_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_1696_), .B(_1692_), .Y(_1697_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(W_151_), .Y(_1698_) );
AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(W_150_), .B(_1083_), .C(_1698_), .Y(_1699_) );
NOR3X1 NOR3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(W_151_), .C(_1087_), .Y(_1700_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1700_), .B(_1699_), .C(_1697_), .Y(_1701_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_1696_), .Y(_1702_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1087_), .B(_788_), .C(W_151_), .Y(_1703_) );
NAND3X1 NAND3X1_201 ( .gnd(gnd), .vdd(vdd), .A(W_150_), .B(_1698_), .C(_1083_), .Y(_1704_) );
NAND3X1 NAND3X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1703_), .B(_1704_), .C(_1702_), .Y(_1705_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .B(_1701_), .Y(_1706_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1706_), .B(_1531_), .Y(_1707_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .Y(_1708_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1708_), .B(_787_), .C(_1095_), .Y(_1709_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_1701_), .B(_1705_), .Y(_1710_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1710_), .B(_1709_), .C(_3610_), .Y(_1711_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(_1707_), .C(W_167_), .Y(_1712_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(W_167_), .Y(_1713_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1530_), .B(_1108_), .C(_1710_), .Y(_1714_) );
AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1706_), .B(_1531_), .C(_3673_), .Y(_1715_) );
NAND3X1 NAND3X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1713_), .B(_1714_), .C(_1715_), .Y(_1716_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1716_), .B(_1712_), .Y(_1717_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .B(_783_), .C(_1457_), .Y(_1718_) );
NAND3X1 NAND3X1_204 ( .gnd(gnd), .vdd(vdd), .A(W_166_), .B(_1463_), .C(_1111_), .Y(_1719_) );
NAND3X1 NAND3X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1718_), .B(_1719_), .C(_1717_), .Y(_1720_) );
NAND3X1 NAND3X1_206 ( .gnd(gnd), .vdd(vdd), .A(W_167_), .B(_1714_), .C(_1715_), .Y(_1721_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(_1707_), .C(_1713_), .Y(_1722_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .B(_1722_), .Y(_1723_) );
AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(W_166_), .B(_1111_), .C(_1463_), .Y(_1724_) );
NOR3X1 NOR3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_1457_), .C(_1115_), .Y(_1725_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .B(_1724_), .C(_1723_), .Y(_1726_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1726_), .B(_1720_), .Y(_1727_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1529_), .B(_1139_), .C(_1727_), .Y(_1728_) );
AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1124_), .B(_1122_), .C(_1529_), .Y(_1729_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_1720_), .B(_1726_), .Y(_1730_) );
AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1729_), .B(_1730_), .C(_3669_), .Y(_1731_) );
NAND3X1 NAND3X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1728_), .C(_1731_), .Y(_1732_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1729_), .B(_1730_), .Y(_1733_) );
AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1118_), .B(_1119_), .C(_654_), .Y(_1734_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1734_), .B(_782_), .C(_1123_), .Y(_1735_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1727_), .B(_1735_), .C(_3617_), .Y(_1736_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .B(_1736_), .C(_1472_), .Y(_1737_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_1732_), .B(_1737_), .Y(_1738_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(W_183_), .Y(_1739_) );
AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(W_182_), .B(_1142_), .C(_1739_), .Y(_1740_) );
AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .B(_1145_), .C(_779_), .Y(_1741_) );
NOR3X1 NOR3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(W_183_), .C(_1741_), .Y(_1742_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1740_), .B(_1742_), .C(_1738_), .Y(_1743_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1732_), .Y(_1744_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1741_), .B(_778_), .C(W_183_), .Y(_1745_) );
NAND3X1 NAND3X1_208 ( .gnd(gnd), .vdd(vdd), .A(W_182_), .B(_1739_), .C(_1142_), .Y(_1746_) );
NAND3X1 NAND3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1745_), .B(_1746_), .C(_1744_), .Y(_1747_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1747_), .B(_1743_), .Y(_1748_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1748_), .B(_1527_), .Y(_1749_) );
AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1150_), .B(_1149_), .C(_673_), .Y(_1750_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1750_), .B(_777_), .C(_1155_), .Y(_1751_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_1743_), .B(_1747_), .Y(_1752_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1752_), .B(_1751_), .C(_3622_), .Y(_1753_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1753_), .B(_1749_), .C(W_199_), .Y(_1754_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(W_199_), .Y(_1755_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1526_), .B(_1172_), .C(_1752_), .Y(_1756_) );
AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1748_), .B(_1527_), .C(_3664_), .Y(_1757_) );
NAND3X1 NAND3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1755_), .B(_1756_), .C(_1757_), .Y(_1758_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1758_), .B(_1754_), .Y(_1759_) );
INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .Y(_1760_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_773_), .C(_1760_), .Y(_1761_) );
NAND3X1 NAND3X1_211 ( .gnd(gnd), .vdd(vdd), .A(W_198_), .B(_1484_), .C(_1175_), .Y(_1762_) );
NAND3X1 NAND3X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1761_), .B(_1762_), .C(_1759_), .Y(_1763_) );
NAND3X1 NAND3X1_213 ( .gnd(gnd), .vdd(vdd), .A(W_199_), .B(_1756_), .C(_1757_), .Y(_1764_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1753_), .B(_1749_), .C(_1755_), .Y(_1765_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1764_), .B(_1765_), .Y(_1766_) );
AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(W_198_), .B(_1175_), .C(_1484_), .Y(_1767_) );
NOR3X1 NOR3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_1760_), .C(_1183_), .Y(_1768_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1768_), .B(_1767_), .C(_1766_), .Y(_1769_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .B(_1763_), .Y(_1770_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1525_), .B(_1770_), .Y(_1771_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_1189_), .Y(_1772_) );
AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1188_), .B(_1190_), .C(_1772_), .Y(_1773_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_1763_), .B(_1769_), .Y(_1774_) );
AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1773_), .B(_1774_), .C(_3660_), .Y(_1775_) );
NAND3X1 NAND3X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1495_), .B(_1771_), .C(_1775_), .Y(_1776_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1773_), .B(_1774_), .Y(_1777_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1770_), .B(_1525_), .C(_3629_), .Y(_1778_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1777_), .B(_1778_), .C(_1496_), .Y(_1780_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_1776_), .B(_1780_), .Y(_1781_) );
INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(W_215_), .Y(_1782_) );
NAND3X1 NAND3X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1209_), .B(_1204_), .C(_1208_), .Y(_1783_) );
AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(W_214_), .B(_1783_), .C(_1782_), .Y(_1784_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(W_215_), .B(_1213_), .Y(_1785_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1785_), .B(_1784_), .C(_1781_), .Y(_1786_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1780_), .B(_1776_), .Y(_1787_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(W_215_), .B(_1213_), .Y(_1788_) );
AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1208_), .B(_1210_), .C(_770_), .Y(_1789_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1782_), .B(_1789_), .Y(_1791_) );
NAND3X1 NAND3X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1787_), .B(_1788_), .C(_1791_), .Y(_1792_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1786_), .B(_1792_), .Y(_1793_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .B(_1793_), .Y(_1794_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1215_), .B(_769_), .C(_1219_), .Y(_1795_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1777_), .B(_1778_), .C(W_215_), .Y(_1796_) );
NAND3X1 NAND3X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1782_), .B(_1771_), .C(_1775_), .Y(_1797_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(W_214_), .B(_1783_), .C(_1797_), .D(_1796_), .Y(_1798_) );
NAND3X1 NAND3X1_218 ( .gnd(gnd), .vdd(vdd), .A(W_215_), .B(_1771_), .C(_1775_), .Y(_1799_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1777_), .B(_1778_), .C(_1782_), .Y(_1800_) );
AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1799_), .B(_1800_), .C(_1213_), .Y(_1802_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1802_), .B(_1798_), .C(_1496_), .Y(_1803_) );
NAND3X1 NAND3X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1799_), .B(_1800_), .C(_1213_), .Y(_1804_) );
NOR3X1 NOR3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1778_), .B(_1782_), .C(_1777_), .Y(_1805_) );
AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1771_), .B(_1775_), .C(W_215_), .Y(_1806_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1805_), .B(_1806_), .C(_1789_), .Y(_1807_) );
NAND3X1 NAND3X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1495_), .B(_1804_), .C(_1807_), .Y(_1808_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(_1808_), .Y(_1809_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1809_), .B(_1795_), .C(_3634_), .Y(_1810_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .B(_1794_), .C(W_231_), .Y(_1811_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(W_231_), .Y(_1813_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1212_), .B(_1239_), .C(_1809_), .Y(_1814_) );
AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .B(_1793_), .C(_3654_), .Y(_1815_) );
NAND3X1 NAND3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1813_), .B(_1814_), .C(_1815_), .Y(_1816_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1816_), .B(_1811_), .Y(_1817_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_765_), .C(_1509_), .Y(_1818_) );
NAND3X1 NAND3X1_222 ( .gnd(gnd), .vdd(vdd), .A(W_230_), .B(_1510_), .C(_1242_), .Y(_1819_) );
NAND3X1 NAND3X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1818_), .B(_1819_), .C(_1817_), .Y(_1820_) );
NAND3X1 NAND3X1_224 ( .gnd(gnd), .vdd(vdd), .A(W_231_), .B(_1814_), .C(_1815_), .Y(_1821_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .B(_1794_), .C(_1813_), .Y(_1822_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1821_), .B(_1822_), .Y(_1824_) );
AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(W_230_), .B(_1242_), .C(_1510_), .Y(_1825_) );
NOR3X1 NOR3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_765_), .B(_1509_), .C(_1246_), .Y(_1826_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1826_), .B(_1825_), .C(_1824_), .Y(_1827_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_1820_), .Y(_1828_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1248_), .B(_1275_), .C(_1828_), .Y(_1829_) );
AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_1254_), .C(_1248_), .Y(_1830_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_1820_), .B(_1827_), .Y(_1831_) );
AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1830_), .B(_1831_), .C(_3641_), .Y(_1832_) );
NAND3X1 NAND3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1522_), .B(_1829_), .C(_1832_), .Y(_1833_) );
INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(_1522_), .Y(_1835_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1830_), .B(_1831_), .Y(_1836_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_3640_), .B(_3638_), .Y(_1837_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1251_), .B(_764_), .C(_1255_), .Y(_1838_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1828_), .B(_1838_), .C(_1837_), .Y(_1839_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1836_), .B(_1839_), .C(_1835_), .Y(_1840_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_1833_), .B(_1840_), .Y(_1841_) );
INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(W_247_), .Y(_1842_) );
AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(W_246_), .B(_1278_), .C(_1842_), .Y(_1843_) );
NOR3X1 NOR3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(W_247_), .C(_1283_), .Y(_1844_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1843_), .B(_1844_), .C(_1841_), .Y(_1846_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1840_), .B(_1833_), .Y(_1847_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(_1280_), .C(W_247_), .Y(_1848_) );
NAND3X1 NAND3X1_226 ( .gnd(gnd), .vdd(vdd), .A(W_246_), .B(_1842_), .C(_1278_), .Y(_1849_) );
NAND3X1 NAND3X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_1849_), .C(_1847_), .Y(_1850_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1850_), .B(_1846_), .Y(_1851_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1851_), .B(_1317_), .Y(_1852_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1852_), .B(_1315_), .Y(_1853_) );
AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1287_), .C(_748_), .Y(_1854_) );
AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1288_), .B(_762_), .C(_1854_), .Y(_1855_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1836_), .B(_1839_), .C(W_247_), .Y(_1857_) );
NAND3X1 NAND3X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(_1829_), .C(_1832_), .Y(_1858_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(W_246_), .B(_1278_), .C(_1858_), .D(_1857_), .Y(_1859_) );
NAND3X1 NAND3X1_229 ( .gnd(gnd), .vdd(vdd), .A(W_247_), .B(_1829_), .C(_1832_), .Y(_1860_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1836_), .B(_1839_), .C(_1842_), .Y(_1861_) );
AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1860_), .B(_1861_), .C(_1279_), .Y(_1862_) );
NOR3X1 NOR3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1835_), .B(_1859_), .C(_1862_), .Y(_1863_) );
NAND3X1 NAND3X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1860_), .B(_1861_), .C(_1279_), .Y(_1864_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_1283_), .Y(_1865_) );
NOR3X1 NOR3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_1842_), .C(_1836_), .Y(_1866_) );
AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1829_), .B(_1832_), .C(W_247_), .Y(_1868_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1866_), .B(_1868_), .C(_1865_), .Y(_1869_) );
AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1864_), .B(_1869_), .C(_1522_), .Y(_1870_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1863_), .B(_1870_), .C(_1855_), .Y(_1871_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1851_), .Y(_1872_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1871_), .B(_1872_), .Y(_1873_) );
NAND3X1 NAND3X1_231 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_1873_), .C(_1312_), .Y(_1874_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1874_), .B(_1853_), .Y(H_7_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_284_), .C(W_248_), .Y(_1875_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(W_248_), .B(_287_), .Y(_1876_) );
INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(_1876_), .Y(_1878_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1875_), .B(_1878_), .Y(H_16_) );
XNOR2X1 XNOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(W_249_), .Y(_1879_) );
XNOR2X1 XNOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1879_), .B(_1878_), .Y(H_17_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_1879_), .Y(_1880_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(W_248_), .B(_287_), .C(_1880_), .Y(_1881_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(W_250_), .Y(_1882_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1882_), .B(_1306_), .Y(_1883_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(W_250_), .B(_1307_), .Y(_1884_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1883_), .B(_1884_), .Y(_1885_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(W_249_), .B(_418_), .C(_1885_), .Y(_1887_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_1887_), .Y(_1888_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(W_249_), .B(_418_), .Y(_1889_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_1889_), .Y(_1890_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1890_), .B(_1885_), .Y(_1891_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1891_), .B(_1888_), .Y(_1892_) );
XNOR2X1 XNOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1892_), .B(_1881_), .Y(H_18_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1891_), .B(_1881_), .C(_1887_), .Y(_1893_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_1883_), .Y(_1894_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(W_251_), .Y(_1895_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1895_), .B(_1522_), .Y(_1897_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(W_251_), .B(_1835_), .Y(_1898_) );
AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1897_), .B(_1898_), .C(_1894_), .Y(_1899_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_1899_), .Y(_1900_) );
NAND3X1 NAND3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1894_), .B(_1897_), .C(_1898_), .Y(_1901_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .B(_1900_), .Y(_1902_) );
XNOR2X1 XNOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .B(_1893_), .Y(H_19_) );
AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .B(_1893_), .C(_1899_), .Y(_1903_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(W_252_), .Y(_1904_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1514_), .B(_1519_), .C(_1517_), .Y(_1905_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1512_), .B(_1509_), .Y(_1907_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1500_), .B(_1319_), .C(_1507_), .Y(_1908_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1321_), .B(_1488_), .C(_1489_), .Y(_1909_) );
INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(_1485_), .Y(_1910_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1481_), .B(_1476_), .C(_1478_), .Y(_1911_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .Y(_1912_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_1465_), .B(_1324_), .Y(_1913_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1462_), .B(_1323_), .C(_1913_), .Y(_1914_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .B(_1326_), .C(_1455_), .Y(_1915_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_1445_), .Y(_1916_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(_1440_), .Y(_1918_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1329_), .B(_1438_), .C(_1918_), .Y(_1919_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1331_), .B(_1423_), .C(_1433_), .Y(_1920_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[92]), .Y(_1921_) );
XNOR2X1 XNOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_2477_), .Y(_1922_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1415_), .B(_1411_), .C(_1413_), .Y(_1923_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1409_), .B(_1406_), .C(_1335_), .Y(_1924_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[76]), .Y(_1925_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_1961_), .Y(_1926_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .Y(_1927_) );
AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1402_), .B(_1403_), .C(_989_), .Y(_1929_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1929_), .B(_1927_), .C(_1404_), .Y(_1930_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[60]), .Y(_1931_) );
XNOR2X1 XNOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_1928_), .Y(_1932_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .Y(_1933_) );
AOI21X1 AOI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1390_), .B(_1338_), .C(_1392_), .Y(_1934_) );
INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(_1934_), .Y(_1935_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[44]), .Y(_1936_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1381_), .B(_1384_), .C(_1378_), .Y(_1937_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[28]), .Y(_1938_) );
XNOR2X1 XNOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_3767_), .B(_1867_), .Y(_1940_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_1940_), .Y(_1941_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1368_), .B(_1369_), .C(_1364_), .Y(_1942_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[12]), .Y(_1943_) );
XNOR2X1 XNOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1834_), .B(_3742_), .Y(_1944_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .Y(_1945_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .Y(_1946_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_1354_), .C(_1946_), .Y(_1947_) );
INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(W_28_), .Y(_1948_) );
XNOR2X1 XNOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(W_0_), .B(W_12_), .Y(_1949_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1949_), .B(W_8_), .Y(_1951_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1948_), .B(_1951_), .Y(_1952_) );
XNOR2X1 XNOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1949_), .B(W_8_), .Y(_1953_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(W_28_), .B(_1953_), .Y(_1954_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1954_), .B(_1952_), .Y(_1955_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(W_27_), .B(W_11_), .C(_1955_), .Y(_1956_) );
XNOR2X1 XNOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1953_), .B(_1948_), .Y(_1957_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(_1957_), .Y(_1958_) );
NAND3X1 NAND3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1947_), .B(_1958_), .C(_1956_), .Y(_1959_) );
AOI21X1 AOI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1958_), .B(_1956_), .C(_1947_), .Y(_1960_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_1960_), .Y(_1962_) );
NAND3X1 NAND3X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1945_), .B(_1959_), .C(_1962_), .Y(_1963_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(_1959_), .Y(_1964_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1964_), .B(_1960_), .C(_1944_), .Y(_1965_) );
NAND3X1 NAND3X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1943_), .B(_1965_), .C(_1963_), .Y(_1966_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1964_), .B(_1960_), .C(_1945_), .Y(_1967_) );
NAND3X1 NAND3X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .B(_1959_), .C(_1962_), .Y(_1968_) );
NAND3X1 NAND3X1_237 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[12]), .B(_1967_), .C(_1968_), .Y(_1969_) );
NAND3X1 NAND3X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .B(_1966_), .C(_1969_), .Y(_1970_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .Y(_1971_) );
NAND3X1 NAND3X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1943_), .B(_1967_), .C(_1968_), .Y(_1973_) );
NAND3X1 NAND3X1_240 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[12]), .B(_1965_), .C(_1963_), .Y(_1974_) );
NAND3X1 NAND3X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_1973_), .C(_1974_), .Y(_1975_) );
NAND3X1 NAND3X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1970_), .B(_1975_), .C(_1942_), .Y(_1976_) );
AOI21X1 AOI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_1344_), .C(_1370_), .Y(_1977_) );
AOI21X1 AOI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1973_), .B(_1974_), .C(_1971_), .Y(_1978_) );
AOI21X1 AOI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .B(_1969_), .C(_1356_), .Y(_1979_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1978_), .B(_1979_), .C(_1977_), .Y(_1980_) );
NAND3X1 NAND3X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1941_), .B(_1976_), .C(_1980_), .Y(_1981_) );
NOR3X1 NOR3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1978_), .B(_1979_), .C(_1977_), .Y(_1982_) );
AOI21X1 AOI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1970_), .B(_1975_), .C(_1942_), .Y(_1984_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1982_), .B(_1984_), .C(_1940_), .Y(_1985_) );
NAND3X1 NAND3X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(_1981_), .C(_1985_), .Y(_1986_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1982_), .B(_1984_), .C(_1941_), .Y(_1987_) );
NAND3X1 NAND3X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1940_), .B(_1976_), .C(_1980_), .Y(_1988_) );
NAND3X1 NAND3X1_246 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[28]), .B(_1988_), .C(_1987_), .Y(_1989_) );
NAND3X1 NAND3X1_247 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .B(_1986_), .C(_1989_), .Y(_1990_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .Y(_1991_) );
NAND3X1 NAND3X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(_1988_), .C(_1987_), .Y(_1992_) );
NAND3X1 NAND3X1_249 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[28]), .B(_1981_), .C(_1985_), .Y(_1993_) );
NAND3X1 NAND3X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1992_), .C(_1993_), .Y(_1995_) );
NAND3X1 NAND3X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_1995_), .C(_1937_), .Y(_1996_) );
AOI21X1 AOI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1376_), .B(_1341_), .C(_1377_), .Y(_1997_) );
AOI21X1 AOI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1992_), .B(_1993_), .C(_1991_), .Y(_1998_) );
AOI21X1 AOI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1986_), .B(_1989_), .C(_1373_), .Y(_1999_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1998_), .B(_1999_), .C(_1997_), .Y(_2000_) );
XNOR2X1 XNOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_1896_), .Y(_2001_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_2001_), .Y(_2002_) );
NAND3X1 NAND3X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_2002_), .C(_2000_), .Y(_2003_) );
NOR3X1 NOR3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1998_), .B(_1997_), .C(_1999_), .Y(_2004_) );
AOI21X1 AOI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_1995_), .C(_1937_), .Y(_2006_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .B(_2006_), .C(_2001_), .Y(_2007_) );
NAND3X1 NAND3X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1936_), .B(_2003_), .C(_2007_), .Y(_2008_) );
NAND3X1 NAND3X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_2001_), .C(_2000_), .Y(_2009_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .B(_2006_), .C(_2002_), .Y(_2010_) );
NAND3X1 NAND3X1_255 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[44]), .B(_2009_), .C(_2010_), .Y(_2011_) );
NAND3X1 NAND3X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1387_), .B(_2008_), .C(_2011_), .Y(_2012_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_1387_), .Y(_2013_) );
NAND3X1 NAND3X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1936_), .B(_2009_), .C(_2010_), .Y(_2014_) );
NAND3X1 NAND3X1_258 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[44]), .B(_2003_), .C(_2007_), .Y(_2015_) );
NAND3X1 NAND3X1_259 ( .gnd(gnd), .vdd(vdd), .A(_2013_), .B(_2014_), .C(_2015_), .Y(_2017_) );
NAND3X1 NAND3X1_260 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(_2017_), .C(_1935_), .Y(_2018_) );
AOI21X1 AOI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_2014_), .B(_2015_), .C(_2013_), .Y(_2019_) );
AOI21X1 AOI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_2008_), .B(_2011_), .C(_1387_), .Y(_2020_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_2019_), .B(_2020_), .C(_1934_), .Y(_2021_) );
NAND3X1 NAND3X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1933_), .B(_2021_), .C(_2018_), .Y(_2022_) );
NOR3X1 NOR3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_2019_), .B(_1934_), .C(_2020_), .Y(_2023_) );
AOI21X1 AOI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(_2017_), .C(_1935_), .Y(_2024_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_2024_), .B(_2023_), .C(_1932_), .Y(_2025_) );
NAND3X1 NAND3X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1931_), .B(_2022_), .C(_2025_), .Y(_2026_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_2024_), .B(_2023_), .C(_1933_), .Y(_2028_) );
NAND3X1 NAND3X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .B(_2021_), .C(_2018_), .Y(_2029_) );
NAND3X1 NAND3X1_264 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[60]), .B(_2029_), .C(_2028_), .Y(_2030_) );
NAND3X1 NAND3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .B(_2026_), .C(_2030_), .Y(_2031_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .Y(_2032_) );
NAND3X1 NAND3X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1931_), .B(_2029_), .C(_2028_), .Y(_2033_) );
NAND3X1 NAND3X1_267 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[60]), .B(_2022_), .C(_2025_), .Y(_2034_) );
NAND3X1 NAND3X1_268 ( .gnd(gnd), .vdd(vdd), .A(_2032_), .B(_2033_), .C(_2034_), .Y(_2035_) );
NAND3X1 NAND3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_2031_), .C(_2035_), .Y(_2036_) );
AOI21X1 AOI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1400_), .B(_1398_), .C(_994_), .Y(_2037_) );
AOI21X1 AOI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1401_), .C(_2037_), .Y(_2039_) );
AOI21X1 AOI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_2033_), .B(_2034_), .C(_2032_), .Y(_2040_) );
AOI21X1 AOI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_2026_), .B(_2030_), .C(_1398_), .Y(_2041_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_2040_), .B(_2041_), .C(_2039_), .Y(_2042_) );
NAND3X1 NAND3X1_270 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .B(_2036_), .C(_2042_), .Y(_2043_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .Y(_2044_) );
NOR3X1 NOR3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_2040_), .B(_2039_), .C(_2041_), .Y(_2045_) );
AOI21X1 AOI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_2031_), .B(_2035_), .C(_1930_), .Y(_2046_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_2045_), .B(_2046_), .C(_2044_), .Y(_2047_) );
NAND3X1 NAND3X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1925_), .B(_2043_), .C(_2047_), .Y(_2048_) );
NAND3X1 NAND3X1_272 ( .gnd(gnd), .vdd(vdd), .A(_2044_), .B(_2036_), .C(_2042_), .Y(_2050_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_2045_), .B(_2046_), .C(_1926_), .Y(_2051_) );
NAND3X1 NAND3X1_273 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[76]), .B(_2050_), .C(_2051_), .Y(_2052_) );
NAND3X1 NAND3X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1924_), .B(_2048_), .C(_2052_), .Y(_2053_) );
INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(_1924_), .Y(_2054_) );
NAND3X1 NAND3X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1925_), .B(_2050_), .C(_2051_), .Y(_2055_) );
NAND3X1 NAND3X1_276 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[76]), .B(_2043_), .C(_2047_), .Y(_2056_) );
NAND3X1 NAND3X1_277 ( .gnd(gnd), .vdd(vdd), .A(_2054_), .B(_2055_), .C(_2056_), .Y(_2057_) );
NAND3X1 NAND3X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1923_), .B(_2053_), .C(_2057_), .Y(_2058_) );
INVX2 INVX2_42 ( .gnd(gnd), .vdd(vdd), .A(_1923_), .Y(_2059_) );
AOI21X1 AOI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_2055_), .B(_2056_), .C(_2054_), .Y(_2061_) );
AOI21X1 AOI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_2048_), .B(_2052_), .C(_1924_), .Y(_2062_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_2061_), .B(_2062_), .C(_2059_), .Y(_2063_) );
NAND3X1 NAND3X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1922_), .B(_2058_), .C(_2063_), .Y(_2064_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(_1922_), .Y(_2065_) );
NAND3X1 NAND3X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1924_), .B(_2055_), .C(_2056_), .Y(_2066_) );
NAND3X1 NAND3X1_281 ( .gnd(gnd), .vdd(vdd), .A(_2054_), .B(_2048_), .C(_2052_), .Y(_2067_) );
AOI21X1 AOI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_2066_), .B(_2067_), .C(_2059_), .Y(_2068_) );
AOI21X1 AOI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_2057_), .C(_1923_), .Y(_2069_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_2068_), .B(_2069_), .C(_2065_), .Y(_2070_) );
NAND3X1 NAND3X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1921_), .B(_2064_), .C(_2070_), .Y(_2072_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_2068_), .B(_2069_), .C(_1922_), .Y(_2073_) );
NAND3X1 NAND3X1_283 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .B(_2058_), .C(_2063_), .Y(_2074_) );
NAND3X1 NAND3X1_284 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[92]), .B(_2074_), .C(_2073_), .Y(_2075_) );
NAND3X1 NAND3X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(_2072_), .C(_2075_), .Y(_2076_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .Y(_2077_) );
NAND3X1 NAND3X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1921_), .B(_2074_), .C(_2073_), .Y(_2078_) );
NAND3X1 NAND3X1_287 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[92]), .B(_2064_), .C(_2070_), .Y(_2079_) );
NAND3X1 NAND3X1_288 ( .gnd(gnd), .vdd(vdd), .A(_2077_), .B(_2078_), .C(_2079_), .Y(_2080_) );
NAND3X1 NAND3X1_289 ( .gnd(gnd), .vdd(vdd), .A(_1920_), .B(_2076_), .C(_2080_), .Y(_2081_) );
AOI21X1 AOI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1432_), .B(_1431_), .C(_1428_), .Y(_2083_) );
AOI21X1 AOI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .B(_2079_), .C(_2077_), .Y(_2084_) );
AOI21X1 AOI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_2072_), .B(_2075_), .C(_1426_), .Y(_2085_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_2084_), .B(_2085_), .C(_2083_), .Y(_2086_) );
NAND3X1 NAND3X1_290 ( .gnd(gnd), .vdd(vdd), .A(_2027_), .B(_2081_), .C(_2086_), .Y(_2087_) );
NOR3X1 NOR3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_2085_), .B(_2083_), .C(_2084_), .Y(_2088_) );
AOI21X1 AOI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_2076_), .B(_2080_), .C(_1920_), .Y(_2089_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_2088_), .B(_2089_), .C(_2444_), .Y(_2090_) );
NAND3X1 NAND3X1_291 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_2087_), .C(_2090_), .Y(_2091_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(W_140_), .B(_2091_), .Y(_2092_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(W_140_), .Y(_2094_) );
NAND3X1 NAND3X1_292 ( .gnd(gnd), .vdd(vdd), .A(_2444_), .B(_2081_), .C(_2086_), .Y(_2095_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_2088_), .B(_2089_), .C(_2027_), .Y(_2096_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_2095_), .B(_2096_), .Y(_2097_) );
NAND3X1 NAND3X1_293 ( .gnd(gnd), .vdd(vdd), .A(_2094_), .B(_116_), .C(_2097_), .Y(_2098_) );
NAND3X1 NAND3X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(_2092_), .C(_2098_), .Y(_2099_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_2094_), .B(_2091_), .Y(_2100_) );
NAND3X1 NAND3X1_295 ( .gnd(gnd), .vdd(vdd), .A(W_140_), .B(_116_), .C(_2097_), .Y(_2101_) );
NAND3X1 NAND3X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1435_), .B(_2100_), .C(_2101_), .Y(_2102_) );
NAND3X1 NAND3X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1919_), .B(_2099_), .C(_2102_), .Y(_2103_) );
INVX2 INVX2_43 ( .gnd(gnd), .vdd(vdd), .A(_1919_), .Y(_2105_) );
AOI21X1 AOI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .B(_2101_), .C(_1435_), .Y(_2106_) );
AOI21X1 AOI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_2092_), .B(_2098_), .C(_1439_), .Y(_2107_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_2107_), .B(_2106_), .C(_2105_), .Y(_2108_) );
NAND3X1 NAND3X1_298 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(_2103_), .C(_2108_), .Y(_2109_) );
NOR3X1 NOR3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_2106_), .B(_2105_), .C(_2107_), .Y(_2110_) );
AOI21X1 AOI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_2099_), .B(_2102_), .C(_1919_), .Y(_2111_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_2110_), .B(_2111_), .C(_2411_), .Y(_2112_) );
NAND3X1 NAND3X1_299 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_2109_), .C(_2112_), .Y(_2113_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(W_156_), .B(_2113_), .Y(_2114_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(W_156_), .Y(_2116_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_2103_), .B(_2108_), .Y(_2117_) );
AOI21X1 AOI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_2411_), .B(_2117_), .C(_143_), .Y(_2118_) );
NAND3X1 NAND3X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2116_), .B(_2109_), .C(_2118_), .Y(_2119_) );
NAND3X1 NAND3X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(_2119_), .C(_2114_), .Y(_2120_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_2116_), .B(_2113_), .Y(_2121_) );
NAND3X1 NAND3X1_302 ( .gnd(gnd), .vdd(vdd), .A(W_156_), .B(_2109_), .C(_2118_), .Y(_2122_) );
NAND3X1 NAND3X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1445_), .B(_2122_), .C(_2121_), .Y(_2123_) );
NAND3X1 NAND3X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2120_), .B(_2123_), .C(_1915_), .Y(_2124_) );
AOI21X1 AOI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1449_), .B(_1454_), .C(_1452_), .Y(_2125_) );
AOI21X1 AOI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_2122_), .B(_2121_), .C(_1445_), .Y(_2127_) );
AOI21X1 AOI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_2119_), .B(_2114_), .C(_1916_), .Y(_2128_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_2128_), .B(_2127_), .C(_2125_), .Y(_2129_) );
AOI21X1 AOI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_2124_), .B(_2129_), .C(_2093_), .Y(_2130_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_2124_), .B(_2129_), .Y(_2131_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_2131_), .B(_2378_), .C(_163_), .Y(_2132_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_2132_), .B(_2130_), .C(W_172_), .Y(_2133_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(W_172_), .Y(_2134_) );
NAND3X1 NAND3X1_305 ( .gnd(gnd), .vdd(vdd), .A(_2378_), .B(_2124_), .C(_2129_), .Y(_2135_) );
NOR3X1 NOR3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_2127_), .B(_2125_), .C(_2128_), .Y(_2136_) );
AOI21X1 AOI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_2120_), .B(_2123_), .C(_1915_), .Y(_2138_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_2136_), .B(_2138_), .C(_2093_), .Y(_2139_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_2135_), .B(_2139_), .Y(_2140_) );
NAND3X1 NAND3X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2134_), .B(_163_), .C(_2140_), .Y(_2141_) );
NAND3X1 NAND3X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1458_), .B(_2133_), .C(_2141_), .Y(_2142_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_2132_), .B(_2130_), .C(_2134_), .Y(_2143_) );
NAND3X1 NAND3X1_308 ( .gnd(gnd), .vdd(vdd), .A(W_172_), .B(_163_), .C(_2140_), .Y(_2144_) );
NAND3X1 NAND3X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_2143_), .C(_2144_), .Y(_2145_) );
NAND3X1 NAND3X1_310 ( .gnd(gnd), .vdd(vdd), .A(_2142_), .B(_2145_), .C(_1914_), .Y(_2146_) );
AOI21X1 AOI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1461_), .B(_1469_), .C(_1466_), .Y(_2147_) );
AOI21X1 AOI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(_2144_), .C(_1464_), .Y(_2149_) );
AOI21X1 AOI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .B(_2141_), .C(_1458_), .Y(_2150_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_2150_), .B(_2149_), .C(_2147_), .Y(_2151_) );
NAND3X1 NAND3X1_311 ( .gnd(gnd), .vdd(vdd), .A(_2126_), .B(_2146_), .C(_2151_), .Y(_2152_) );
NOR3X1 NOR3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_2149_), .B(_2147_), .C(_2150_), .Y(_2153_) );
AOI21X1 AOI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_2142_), .B(_2145_), .C(_1914_), .Y(_2154_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_2153_), .B(_2154_), .C(_2356_), .Y(_2155_) );
NAND3X1 NAND3X1_312 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_2152_), .C(_2155_), .Y(_2156_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(W_188_), .B(_2156_), .Y(_2157_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(W_188_), .Y(_2158_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_2146_), .B(_2151_), .Y(_2160_) );
AOI21X1 AOI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_2356_), .B(_2160_), .C(_191_), .Y(_2161_) );
NAND3X1 NAND3X1_313 ( .gnd(gnd), .vdd(vdd), .A(_2158_), .B(_2152_), .C(_2161_), .Y(_2162_) );
NAND3X1 NAND3X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(_2162_), .C(_2157_), .Y(_2163_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_2158_), .B(_2156_), .Y(_2164_) );
NAND3X1 NAND3X1_315 ( .gnd(gnd), .vdd(vdd), .A(W_188_), .B(_2152_), .C(_2161_), .Y(_2165_) );
NAND3X1 NAND3X1_316 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(_2165_), .C(_2164_), .Y(_2166_) );
NAND3X1 NAND3X1_317 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(_2166_), .C(_1911_), .Y(_2167_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(_1478_), .Y(_2168_) );
AOI21X1 AOI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1322_), .B(_1477_), .C(_2168_), .Y(_2169_) );
AOI21X1 AOI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_2165_), .B(_2164_), .C(_1473_), .Y(_2171_) );
AOI21X1 AOI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_2162_), .B(_2157_), .C(_1912_), .Y(_2172_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_2171_), .B(_2172_), .C(_2169_), .Y(_2173_) );
NAND3X1 NAND3X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2159_), .B(_2167_), .C(_2173_), .Y(_2174_) );
NOR3X1 NOR3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_2171_), .B(_2172_), .C(_2169_), .Y(_2175_) );
AOI21X1 AOI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(_2166_), .C(_1911_), .Y(_2176_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_2175_), .B(_2176_), .C(_2334_), .Y(_2177_) );
NAND3X1 NAND3X1_319 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_2174_), .C(_2177_), .Y(_2178_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(W_204_), .B(_2178_), .Y(_2179_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(W_204_), .Y(_2180_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_2167_), .B(_2173_), .Y(_2182_) );
AOI21X1 AOI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_2334_), .B(_2182_), .C(_217_), .Y(_2183_) );
NAND3X1 NAND3X1_320 ( .gnd(gnd), .vdd(vdd), .A(_2180_), .B(_2174_), .C(_2183_), .Y(_2184_) );
NAND3X1 NAND3X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1910_), .B(_2184_), .C(_2179_), .Y(_2185_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_2180_), .B(_2178_), .Y(_2186_) );
NAND3X1 NAND3X1_322 ( .gnd(gnd), .vdd(vdd), .A(W_204_), .B(_2174_), .C(_2183_), .Y(_2187_) );
NAND3X1 NAND3X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1485_), .B(_2187_), .C(_2186_), .Y(_2188_) );
NAND3X1 NAND3X1_324 ( .gnd(gnd), .vdd(vdd), .A(_2185_), .B(_1909_), .C(_2188_), .Y(_2189_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1227_), .B(_399_), .C(_1232_), .Y(_2190_) );
AOI21X1 AOI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_2190_), .B(_1492_), .C(_1490_), .Y(_2191_) );
AOI21X1 AOI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_2187_), .B(_2186_), .C(_1485_), .Y(_2193_) );
AOI21X1 AOI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_2184_), .B(_2179_), .C(_1910_), .Y(_2194_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_2193_), .B(_2194_), .C(_2191_), .Y(_2195_) );
NAND3X1 NAND3X1_325 ( .gnd(gnd), .vdd(vdd), .A(_2192_), .B(_2189_), .C(_2195_), .Y(_2196_) );
NAND3X1 NAND3X1_326 ( .gnd(gnd), .vdd(vdd), .A(_1485_), .B(_2184_), .C(_2179_), .Y(_2197_) );
NAND3X1 NAND3X1_327 ( .gnd(gnd), .vdd(vdd), .A(_1910_), .B(_2187_), .C(_2186_), .Y(_2198_) );
AOI21X1 AOI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_2197_), .B(_2198_), .C(_2191_), .Y(_2199_) );
AOI21X1 AOI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_2185_), .B(_2188_), .C(_1909_), .Y(_2200_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_2199_), .B(_2200_), .C(_2312_), .Y(_2201_) );
NAND3X1 NAND3X1_328 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_2196_), .C(_2201_), .Y(_2202_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(W_220_), .B(_2202_), .Y(_2204_) );
INVX2 INVX2_44 ( .gnd(gnd), .vdd(vdd), .A(W_220_), .Y(_2205_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_2201_), .B(_236_), .Y(_2206_) );
NAND3X1 NAND3X1_329 ( .gnd(gnd), .vdd(vdd), .A(_2205_), .B(_2196_), .C(_2206_), .Y(_2207_) );
NAND3X1 NAND3X1_330 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_2204_), .C(_2207_), .Y(_2208_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_2205_), .B(_2202_), .Y(_2209_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_2202_), .B(_2205_), .Y(_2210_) );
NAND3X1 NAND3X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1497_), .B(_2209_), .C(_2210_), .Y(_2211_) );
NAND3X1 NAND3X1_332 ( .gnd(gnd), .vdd(vdd), .A(_2208_), .B(_2211_), .C(_1908_), .Y(_2212_) );
AOI21X1 AOI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .B(_1505_), .C(_1503_), .Y(_2213_) );
AOI21X1 AOI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_2209_), .B(_2210_), .C(_1497_), .Y(_2215_) );
AOI21X1 AOI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_2204_), .B(_2207_), .C(_1502_), .Y(_2216_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_2215_), .B(_2216_), .C(_2213_), .Y(_2217_) );
NAND3X1 NAND3X1_333 ( .gnd(gnd), .vdd(vdd), .A(_2225_), .B(_2212_), .C(_2217_), .Y(_2218_) );
NAND3X1 NAND3X1_334 ( .gnd(gnd), .vdd(vdd), .A(_1497_), .B(_2204_), .C(_2207_), .Y(_2219_) );
NAND3X1 NAND3X1_335 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_2209_), .C(_2210_), .Y(_2220_) );
AOI21X1 AOI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_2219_), .B(_2220_), .C(_2213_), .Y(_2221_) );
AOI21X1 AOI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_2208_), .B(_2211_), .C(_1908_), .Y(_2222_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_2222_), .B(_2221_), .C(_2290_), .Y(_2223_) );
NAND3X1 NAND3X1_336 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_2218_), .C(_2223_), .Y(_2224_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(W_236_), .B(_2224_), .Y(_2226_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(W_236_), .Y(_2227_) );
NAND3X1 NAND3X1_337 ( .gnd(gnd), .vdd(vdd), .A(_2290_), .B(_2212_), .C(_2217_), .Y(_2228_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_2222_), .B(_2221_), .C(_2225_), .Y(_2229_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_2228_), .B(_2229_), .Y(_2230_) );
NAND3X1 NAND3X1_338 ( .gnd(gnd), .vdd(vdd), .A(_2227_), .B(_261_), .C(_2230_), .Y(_2231_) );
NAND3X1 NAND3X1_339 ( .gnd(gnd), .vdd(vdd), .A(_1907_), .B(_2226_), .C(_2231_), .Y(_2232_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_2227_), .B(_2224_), .Y(_2233_) );
NAND3X1 NAND3X1_340 ( .gnd(gnd), .vdd(vdd), .A(W_236_), .B(_261_), .C(_2230_), .Y(_2234_) );
NAND3X1 NAND3X1_341 ( .gnd(gnd), .vdd(vdd), .A(_1511_), .B(_2233_), .C(_2234_), .Y(_2235_) );
NAND3X1 NAND3X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2232_), .B(_2235_), .C(_1905_), .Y(_2237_) );
AOI21X1 AOI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1318_), .B(_1515_), .C(_1520_), .Y(_2238_) );
AOI21X1 AOI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_2233_), .B(_2234_), .C(_1511_), .Y(_2239_) );
AOI21X1 AOI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_2226_), .B(_2231_), .C(_1907_), .Y(_2240_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_2239_), .B(_2240_), .C(_2238_), .Y(_2241_) );
AOI21X1 AOI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_2241_), .B(_2237_), .C(_2257_), .Y(_2242_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_2241_), .B(_2237_), .Y(_2243_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_2243_), .B(_2268_), .C(_286_), .Y(_2244_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_2244_), .B(_2242_), .C(_1904_), .Y(_2245_) );
NOR3X1 NOR3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_2239_), .B(_2240_), .C(_2238_), .Y(_2246_) );
AOI21X1 AOI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_2232_), .B(_2235_), .C(_1905_), .Y(_2248_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_2246_), .B(_2248_), .C(_2257_), .Y(_2249_) );
NAND3X1 NAND3X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2268_), .B(_2241_), .C(_2237_), .Y(_2250_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_2250_), .B(_2249_), .Y(_2251_) );
NAND3X1 NAND3X1_344 ( .gnd(gnd), .vdd(vdd), .A(W_252_), .B(_286_), .C(_2251_), .Y(_2252_) );
NAND3X1 NAND3X1_345 ( .gnd(gnd), .vdd(vdd), .A(_1897_), .B(_2245_), .C(_2252_), .Y(_2253_) );
AOI21X1 AOI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_2245_), .B(_2252_), .C(_1897_), .Y(_2254_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_2254_), .Y(_2255_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_2253_), .B(_2255_), .Y(_2256_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_2256_), .B(_1903_), .Y(H_20_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_2254_), .B(_1903_), .C(_2253_), .Y(_2258_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_2251_), .Y(_2259_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(W_252_), .B(_2259_), .Y(_2260_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(W_253_), .Y(_2261_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_2238_), .B(_2240_), .C(_2232_), .Y(_2262_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(W_237_), .Y(_2263_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_2216_), .B(_2213_), .C(_2208_), .Y(_2264_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(W_221_), .Y(_2265_) );
AOI21X1 AOI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_2188_), .B(_1909_), .C(_2193_), .Y(_2266_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(_2179_), .Y(_2267_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(W_205_), .Y(_2269_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_2169_), .B(_2172_), .C(_2163_), .Y(_2270_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(W_189_), .Y(_2271_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_2150_), .B(_2147_), .C(_2142_), .Y(_2272_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(W_173_), .Y(_2273_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_3206_), .Y(_2274_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_2128_), .B(_2125_), .C(_2120_), .Y(_2275_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(W_157_), .Y(_2276_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(_3198_), .Y(_2277_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_2107_), .B(_2105_), .C(_2099_), .Y(_2278_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(W_141_), .Y(_2280_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_2085_), .B(_2083_), .C(_2076_), .Y(_2281_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_2059_), .B(_2062_), .C(_2053_), .Y(_2282_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_2041_), .B(_2039_), .C(_2031_), .Y(_2283_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_2020_), .B(_1934_), .C(_2012_), .Y(_2284_) );
AOI21X1 AOI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1995_), .B(_1937_), .C(_1998_), .Y(_2285_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[29]), .Y(_2286_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1977_), .B(_1979_), .C(_1970_), .Y(_2287_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(_1957_), .Y(_2288_) );
AOI21X1 AOI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1947_), .B(_1958_), .C(_2288_), .Y(_2289_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(_1952_), .Y(_2291_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(W_29_), .Y(_2292_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(W_12_), .B(W_13_), .Y(_2293_) );
XNOR2X1 XNOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_314_), .Y(_2294_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .B(_2294_), .Y(_2295_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .Y(_2296_) );
XNOR2X1 XNOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(W_9_), .Y(_2297_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_2296_), .B(_2297_), .Y(_2298_) );
AOI21X1 AOI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_2295_), .B(_2298_), .C(_2292_), .Y(_2299_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_2296_), .B(_2294_), .Y(_2300_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .B(_2297_), .Y(_2302_) );
AOI21X1 AOI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_2300_), .B(_2302_), .C(W_29_), .Y(_2303_) );
NOR3X1 NOR3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_2299_), .B(_2291_), .C(_2303_), .Y(_2304_) );
NAND3X1 NAND3X1_346 ( .gnd(gnd), .vdd(vdd), .A(W_29_), .B(_2300_), .C(_2302_), .Y(_2305_) );
NAND3X1 NAND3X1_347 ( .gnd(gnd), .vdd(vdd), .A(_2292_), .B(_2295_), .C(_2298_), .Y(_2306_) );
AOI21X1 AOI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_2305_), .B(_2306_), .C(_1952_), .Y(_2307_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_2304_), .B(_2307_), .C(_2289_), .Y(_2308_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(_1947_), .Y(_2309_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1351_), .B(_1955_), .Y(_2310_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_2309_), .B(_2310_), .C(_1956_), .Y(_2311_) );
NAND3X1 NAND3X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1952_), .B(_2305_), .C(_2306_), .Y(_2313_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_2299_), .B(_2303_), .C(_2291_), .Y(_2314_) );
NAND3X1 NAND3X1_349 ( .gnd(gnd), .vdd(vdd), .A(_2313_), .B(_2314_), .C(_2311_), .Y(_2315_) );
XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_2751_), .B(_321_), .Y(_2316_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(_2316_), .Y(_2317_) );
NAND3X1 NAND3X1_350 ( .gnd(gnd), .vdd(vdd), .A(_2308_), .B(_2317_), .C(_2315_), .Y(_2318_) );
AOI21X1 AOI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_2313_), .B(_2314_), .C(_2311_), .Y(_2319_) );
NOR3X1 NOR3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_2289_), .B(_2307_), .C(_2304_), .Y(_2320_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_2320_), .B(_2319_), .C(_2316_), .Y(_2321_) );
NAND3X1 NAND3X1_351 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[13]), .B(_2318_), .C(_2321_), .Y(_2322_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[13]), .Y(_2324_) );
NOR3X1 NOR3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_2319_), .B(_2316_), .C(_2320_), .Y(_2325_) );
AOI21X1 AOI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_2308_), .B(_2315_), .C(_2317_), .Y(_2326_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_2325_), .B(_2326_), .C(_2324_), .Y(_2327_) );
NAND3X1 NAND3X1_352 ( .gnd(gnd), .vdd(vdd), .A(_1973_), .B(_2322_), .C(_2327_), .Y(_2328_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(_1973_), .Y(_2329_) );
NOR3X1 NOR3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_2324_), .B(_2326_), .C(_2325_), .Y(_2330_) );
AOI21X1 AOI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_2318_), .B(_2321_), .C(bloque_datos[13]), .Y(_2331_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_2330_), .B(_2331_), .C(_2329_), .Y(_2332_) );
NAND3X1 NAND3X1_353 ( .gnd(gnd), .vdd(vdd), .A(_2328_), .B(_2287_), .C(_2332_), .Y(_2333_) );
AOI21X1 AOI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1975_), .B(_1942_), .C(_1978_), .Y(_2335_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_2330_), .B(_2331_), .C(_1973_), .Y(_2336_) );
NAND3X1 NAND3X1_354 ( .gnd(gnd), .vdd(vdd), .A(_2329_), .B(_2322_), .C(_2327_), .Y(_2337_) );
NAND3X1 NAND3X1_355 ( .gnd(gnd), .vdd(vdd), .A(_2337_), .B(_2335_), .C(_2336_), .Y(_2338_) );
XNOR2X1 XNOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_496_), .Y(_2339_) );
NAND3X1 NAND3X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .B(_2338_), .C(_2333_), .Y(_2340_) );
AOI21X1 AOI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_2337_), .B(_2336_), .C(_2335_), .Y(_2341_) );
AOI21X1 AOI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_2328_), .B(_2332_), .C(_2287_), .Y(_2342_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .Y(_2343_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_2341_), .B(_2342_), .C(_2343_), .Y(_2344_) );
AOI21X1 AOI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_2340_), .B(_2344_), .C(_2286_), .Y(_2346_) );
NAND3X1 NAND3X1_357 ( .gnd(gnd), .vdd(vdd), .A(_2343_), .B(_2338_), .C(_2333_), .Y(_2347_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_2341_), .B(_2342_), .C(_2339_), .Y(_2348_) );
AOI21X1 AOI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_2347_), .B(_2348_), .C(bloque_datos[29]), .Y(_2349_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_2346_), .B(_2349_), .C(_1992_), .Y(_2350_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(_1992_), .Y(_2351_) );
NAND3X1 NAND3X1_358 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[29]), .B(_2347_), .C(_2348_), .Y(_2352_) );
NAND3X1 NAND3X1_359 ( .gnd(gnd), .vdd(vdd), .A(_2286_), .B(_2340_), .C(_2344_), .Y(_2353_) );
NAND3X1 NAND3X1_360 ( .gnd(gnd), .vdd(vdd), .A(_2351_), .B(_2352_), .C(_2353_), .Y(_2354_) );
AOI21X1 AOI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_2354_), .B(_2350_), .C(_2285_), .Y(_2355_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1999_), .B(_1997_), .C(_1990_), .Y(_2357_) );
NAND3X1 NAND3X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1992_), .B(_2352_), .C(_2353_), .Y(_2358_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_2346_), .B(_2349_), .C(_2351_), .Y(_2359_) );
AOI21X1 AOI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_2358_), .B(_2359_), .C(_2357_), .Y(_2360_) );
XNOR2X1 XNOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_2905_), .Y(_2361_) );
NOR3X1 NOR3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_2355_), .B(_2361_), .C(_2360_), .Y(_2362_) );
NAND3X1 NAND3X1_362 ( .gnd(gnd), .vdd(vdd), .A(_2358_), .B(_2357_), .C(_2359_), .Y(_2363_) );
NAND3X1 NAND3X1_363 ( .gnd(gnd), .vdd(vdd), .A(_2354_), .B(_2285_), .C(_2350_), .Y(_2364_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(_2361_), .Y(_2365_) );
AOI21X1 AOI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_2363_), .B(_2364_), .C(_2365_), .Y(_2366_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_2362_), .B(_2366_), .C(bloque_datos[45]), .Y(_2368_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[45]), .Y(_2369_) );
NAND3X1 NAND3X1_364 ( .gnd(gnd), .vdd(vdd), .A(_2365_), .B(_2363_), .C(_2364_), .Y(_2370_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_2360_), .B(_2355_), .C(_2361_), .Y(_2371_) );
NAND3X1 NAND3X1_365 ( .gnd(gnd), .vdd(vdd), .A(_2369_), .B(_2370_), .C(_2371_), .Y(_2372_) );
NAND3X1 NAND3X1_366 ( .gnd(gnd), .vdd(vdd), .A(_2014_), .B(_2372_), .C(_2368_), .Y(_2373_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(_2014_), .Y(_2374_) );
AOI21X1 AOI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_2370_), .B(_2371_), .C(_2369_), .Y(_2375_) );
NOR3X1 NOR3X1_45 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[45]), .B(_2366_), .C(_2362_), .Y(_2376_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_2376_), .B(_2375_), .C(_2374_), .Y(_2377_) );
NAND3X1 NAND3X1_367 ( .gnd(gnd), .vdd(vdd), .A(_2373_), .B(_2284_), .C(_2377_), .Y(_2379_) );
AOI21X1 AOI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_2017_), .B(_1935_), .C(_2019_), .Y(_2380_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_2376_), .B(_2375_), .C(_2014_), .Y(_2381_) );
NAND3X1 NAND3X1_368 ( .gnd(gnd), .vdd(vdd), .A(_2374_), .B(_2372_), .C(_2368_), .Y(_2382_) );
NAND3X1 NAND3X1_369 ( .gnd(gnd), .vdd(vdd), .A(_2381_), .B(_2382_), .C(_2380_), .Y(_2383_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_2949_), .B(_2959_), .Y(_2384_) );
XNOR2X1 XNOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_2384_), .Y(_2385_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(_2385_), .Y(_2386_) );
NAND3X1 NAND3X1_370 ( .gnd(gnd), .vdd(vdd), .A(_2379_), .B(_2386_), .C(_2383_), .Y(_2387_) );
AOI21X1 AOI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_2382_), .B(_2381_), .C(_2380_), .Y(_2388_) );
AOI21X1 AOI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_2373_), .B(_2377_), .C(_2284_), .Y(_2390_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_2388_), .B(_2390_), .C(_2385_), .Y(_2391_) );
NAND3X1 NAND3X1_371 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[61]), .B(_2387_), .C(_2391_), .Y(_2392_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[61]), .Y(_2393_) );
NAND3X1 NAND3X1_372 ( .gnd(gnd), .vdd(vdd), .A(_2379_), .B(_2385_), .C(_2383_), .Y(_2394_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_2388_), .B(_2390_), .C(_2386_), .Y(_2395_) );
NAND3X1 NAND3X1_373 ( .gnd(gnd), .vdd(vdd), .A(_2393_), .B(_2394_), .C(_2395_), .Y(_2396_) );
NAND3X1 NAND3X1_374 ( .gnd(gnd), .vdd(vdd), .A(_2033_), .B(_2392_), .C(_2396_), .Y(_2397_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(_2033_), .Y(_2398_) );
AOI21X1 AOI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_2394_), .B(_2395_), .C(_2393_), .Y(_2399_) );
AOI21X1 AOI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_2387_), .B(_2391_), .C(bloque_datos[61]), .Y(_2401_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .B(_2401_), .C(_2398_), .Y(_2402_) );
NAND3X1 NAND3X1_375 ( .gnd(gnd), .vdd(vdd), .A(_2283_), .B(_2397_), .C(_2402_), .Y(_2403_) );
AOI21X1 AOI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_2035_), .C(_2040_), .Y(_2404_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .B(_2401_), .C(_2033_), .Y(_2405_) );
NAND3X1 NAND3X1_376 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .B(_2392_), .C(_2396_), .Y(_2406_) );
NAND3X1 NAND3X1_377 ( .gnd(gnd), .vdd(vdd), .A(_2404_), .B(_2406_), .C(_2405_), .Y(_2407_) );
XNOR2X1 XNOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_3080_), .Y(_2408_) );
NAND3X1 NAND3X1_378 ( .gnd(gnd), .vdd(vdd), .A(_2408_), .B(_2403_), .C(_2407_), .Y(_2409_) );
AOI21X1 AOI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_2406_), .B(_2405_), .C(_2404_), .Y(_2410_) );
AOI21X1 AOI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_2397_), .B(_2402_), .C(_2283_), .Y(_2412_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(_2408_), .Y(_2413_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_2410_), .B(_2412_), .C(_2413_), .Y(_2414_) );
NAND3X1 NAND3X1_379 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[77]), .B(_2409_), .C(_2414_), .Y(_2415_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[77]), .Y(_2416_) );
NAND3X1 NAND3X1_380 ( .gnd(gnd), .vdd(vdd), .A(_2413_), .B(_2403_), .C(_2407_), .Y(_2417_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_2410_), .B(_2412_), .C(_2408_), .Y(_2418_) );
NAND3X1 NAND3X1_381 ( .gnd(gnd), .vdd(vdd), .A(_2416_), .B(_2417_), .C(_2418_), .Y(_2419_) );
NAND3X1 NAND3X1_382 ( .gnd(gnd), .vdd(vdd), .A(_2055_), .B(_2415_), .C(_2419_), .Y(_2420_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(_2055_), .Y(_2421_) );
AOI21X1 AOI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_2417_), .B(_2418_), .C(_2416_), .Y(_2423_) );
AOI21X1 AOI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_2409_), .B(_2414_), .C(bloque_datos[77]), .Y(_2424_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_2423_), .B(_2424_), .C(_2421_), .Y(_2425_) );
NAND3X1 NAND3X1_383 ( .gnd(gnd), .vdd(vdd), .A(_2420_), .B(_2425_), .C(_2282_), .Y(_2426_) );
AOI21X1 AOI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1923_), .B(_2057_), .C(_2061_), .Y(_2427_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_2423_), .B(_2424_), .C(_2055_), .Y(_2428_) );
NAND3X1 NAND3X1_384 ( .gnd(gnd), .vdd(vdd), .A(_2421_), .B(_2415_), .C(_2419_), .Y(_2429_) );
NAND3X1 NAND3X1_385 ( .gnd(gnd), .vdd(vdd), .A(_2429_), .B(_2427_), .C(_2428_), .Y(_2430_) );
XNOR2X1 XNOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_3146_), .Y(_2431_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(_2431_), .Y(_2432_) );
NAND3X1 NAND3X1_386 ( .gnd(gnd), .vdd(vdd), .A(_2432_), .B(_2430_), .C(_2426_), .Y(_2434_) );
AOI21X1 AOI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_2429_), .B(_2428_), .C(_2427_), .Y(_2435_) );
AOI21X1 AOI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_2420_), .B(_2425_), .C(_2282_), .Y(_2436_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_2435_), .B(_2436_), .C(_2431_), .Y(_2437_) );
NAND3X1 NAND3X1_387 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[93]), .B(_2434_), .C(_2437_), .Y(_2438_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[93]), .Y(_2439_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_2435_), .B(_2436_), .C(_2432_), .Y(_2440_) );
NAND3X1 NAND3X1_388 ( .gnd(gnd), .vdd(vdd), .A(_2431_), .B(_2430_), .C(_2426_), .Y(_2441_) );
NAND3X1 NAND3X1_389 ( .gnd(gnd), .vdd(vdd), .A(_2439_), .B(_2441_), .C(_2440_), .Y(_2442_) );
NAND3X1 NAND3X1_390 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .B(_2438_), .C(_2442_), .Y(_2443_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .Y(_2445_) );
AOI21X1 AOI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_2441_), .B(_2440_), .C(_2439_), .Y(_2446_) );
AOI21X1 AOI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_2434_), .B(_2437_), .C(bloque_datos[93]), .Y(_2447_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_2446_), .B(_2447_), .C(_2445_), .Y(_2448_) );
NAND3X1 NAND3X1_391 ( .gnd(gnd), .vdd(vdd), .A(_2443_), .B(_2281_), .C(_2448_), .Y(_2449_) );
AOI21X1 AOI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1920_), .B(_2080_), .C(_2084_), .Y(_2450_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_2446_), .B(_2447_), .C(_2078_), .Y(_2451_) );
NAND3X1 NAND3X1_392 ( .gnd(gnd), .vdd(vdd), .A(_2445_), .B(_2438_), .C(_2442_), .Y(_2452_) );
NAND3X1 NAND3X1_393 ( .gnd(gnd), .vdd(vdd), .A(_2450_), .B(_2452_), .C(_2451_), .Y(_2453_) );
AOI21X1 AOI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_2449_), .B(_2453_), .C(_3190_), .Y(_2454_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(_2454_), .Y(_2456_) );
NAND3X1 NAND3X1_394 ( .gnd(gnd), .vdd(vdd), .A(_3190_), .B(_2449_), .C(_2453_), .Y(_2457_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_2457_), .B(_360_), .Y(_2458_) );
NAND3X1 NAND3X1_395 ( .gnd(gnd), .vdd(vdd), .A(_2280_), .B(_2456_), .C(_2458_), .Y(_2459_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_2457_), .Y(_2460_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_2460_), .B(_2454_), .C(W_141_), .Y(_2461_) );
NAND3X1 NAND3X1_396 ( .gnd(gnd), .vdd(vdd), .A(_2092_), .B(_2461_), .C(_2459_), .Y(_2462_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(_2092_), .Y(_2463_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_2460_), .B(_2454_), .C(_2280_), .Y(_2464_) );
NAND3X1 NAND3X1_397 ( .gnd(gnd), .vdd(vdd), .A(W_141_), .B(_2456_), .C(_2458_), .Y(_2465_) );
NAND3X1 NAND3X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2463_), .B(_2464_), .C(_2465_), .Y(_2467_) );
NAND3X1 NAND3X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2462_), .B(_2467_), .C(_2278_), .Y(_2468_) );
AOI21X1 AOI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1919_), .B(_2102_), .C(_2106_), .Y(_2469_) );
AOI21X1 AOI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_2464_), .B(_2465_), .C(_2463_), .Y(_2470_) );
AOI21X1 AOI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_2461_), .B(_2459_), .C(_2092_), .Y(_2471_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .B(_2471_), .C(_2469_), .Y(_2472_) );
NAND3X1 NAND3X1_400 ( .gnd(gnd), .vdd(vdd), .A(_2277_), .B(_2468_), .C(_2472_), .Y(_2473_) );
NOR3X1 NOR3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .B(_2469_), .C(_2471_), .Y(_2474_) );
AOI21X1 AOI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_2462_), .B(_2467_), .C(_2278_), .Y(_2475_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_2474_), .B(_2475_), .C(_3198_), .Y(_2476_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .B(_2476_), .Y(_2478_) );
NAND3X1 NAND3X1_401 ( .gnd(gnd), .vdd(vdd), .A(_2276_), .B(_369_), .C(_2478_), .Y(_2479_) );
NAND3X1 NAND3X1_402 ( .gnd(gnd), .vdd(vdd), .A(_3198_), .B(_2468_), .C(_2472_), .Y(_2480_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_2474_), .B(_2475_), .C(_2277_), .Y(_2481_) );
NAND3X1 NAND3X1_403 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_2480_), .C(_2481_), .Y(_2482_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(W_157_), .B(_2482_), .Y(_2483_) );
NAND3X1 NAND3X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2114_), .B(_2479_), .C(_2483_), .Y(_2484_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(_2114_), .Y(_2485_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_2276_), .B(_2482_), .Y(_2486_) );
NAND3X1 NAND3X1_405 ( .gnd(gnd), .vdd(vdd), .A(W_157_), .B(_369_), .C(_2478_), .Y(_2487_) );
NAND3X1 NAND3X1_406 ( .gnd(gnd), .vdd(vdd), .A(_2485_), .B(_2486_), .C(_2487_), .Y(_2489_) );
NAND3X1 NAND3X1_407 ( .gnd(gnd), .vdd(vdd), .A(_2275_), .B(_2484_), .C(_2489_), .Y(_2490_) );
AOI21X1 AOI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_2123_), .B(_1915_), .C(_2127_), .Y(_2491_) );
AOI21X1 AOI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_2486_), .B(_2487_), .C(_2485_), .Y(_2492_) );
AOI21X1 AOI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_2479_), .B(_2483_), .C(_2114_), .Y(_2493_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_2492_), .B(_2493_), .C(_2491_), .Y(_2494_) );
NAND3X1 NAND3X1_408 ( .gnd(gnd), .vdd(vdd), .A(_2274_), .B(_2490_), .C(_2494_), .Y(_2495_) );
NOR3X1 NOR3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_2492_), .B(_2491_), .C(_2493_), .Y(_2496_) );
AOI21X1 AOI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .B(_2489_), .C(_2275_), .Y(_2497_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_2496_), .B(_2497_), .C(_3206_), .Y(_2498_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_2495_), .B(_2498_), .Y(_2500_) );
NAND3X1 NAND3X1_409 ( .gnd(gnd), .vdd(vdd), .A(_2273_), .B(_378_), .C(_2500_), .Y(_2501_) );
NAND3X1 NAND3X1_410 ( .gnd(gnd), .vdd(vdd), .A(_3206_), .B(_2490_), .C(_2494_), .Y(_2502_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_2496_), .B(_2497_), .C(_2274_), .Y(_2503_) );
NAND3X1 NAND3X1_411 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_2502_), .C(_2503_), .Y(_2504_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(W_173_), .B(_2504_), .Y(_2505_) );
NAND3X1 NAND3X1_412 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .B(_2501_), .C(_2505_), .Y(_2506_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .Y(_2507_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_2273_), .B(_2504_), .Y(_2508_) );
NAND3X1 NAND3X1_413 ( .gnd(gnd), .vdd(vdd), .A(W_173_), .B(_378_), .C(_2500_), .Y(_2509_) );
NAND3X1 NAND3X1_414 ( .gnd(gnd), .vdd(vdd), .A(_2507_), .B(_2508_), .C(_2509_), .Y(_2511_) );
NAND3X1 NAND3X1_415 ( .gnd(gnd), .vdd(vdd), .A(_2272_), .B(_2506_), .C(_2511_), .Y(_2512_) );
AOI21X1 AOI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_2145_), .B(_1914_), .C(_2149_), .Y(_2513_) );
AOI21X1 AOI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_2508_), .B(_2509_), .C(_2507_), .Y(_2514_) );
AOI21X1 AOI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .B(_2505_), .C(_2133_), .Y(_2515_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_2514_), .B(_2515_), .C(_2513_), .Y(_2516_) );
NAND3X1 NAND3X1_416 ( .gnd(gnd), .vdd(vdd), .A(_3216_), .B(_2512_), .C(_2516_), .Y(_2517_) );
NOR3X1 NOR3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_2514_), .B(_2513_), .C(_2515_), .Y(_2518_) );
AOI21X1 AOI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_2506_), .B(_2511_), .C(_2272_), .Y(_2519_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_2518_), .B(_2519_), .C(_3214_), .Y(_2520_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_2517_), .B(_2520_), .Y(_2522_) );
NAND3X1 NAND3X1_417 ( .gnd(gnd), .vdd(vdd), .A(_2271_), .B(_386_), .C(_2522_), .Y(_2523_) );
NAND3X1 NAND3X1_418 ( .gnd(gnd), .vdd(vdd), .A(_3214_), .B(_2512_), .C(_2516_), .Y(_2524_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_2518_), .B(_2519_), .C(_3216_), .Y(_2525_) );
NAND3X1 NAND3X1_419 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_2524_), .C(_2525_), .Y(_2526_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(W_189_), .B(_2526_), .Y(_2527_) );
NAND3X1 NAND3X1_420 ( .gnd(gnd), .vdd(vdd), .A(_2157_), .B(_2523_), .C(_2527_), .Y(_2528_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(_2157_), .Y(_2529_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_2271_), .B(_2526_), .Y(_2530_) );
NAND3X1 NAND3X1_421 ( .gnd(gnd), .vdd(vdd), .A(W_189_), .B(_386_), .C(_2522_), .Y(_2531_) );
NAND3X1 NAND3X1_422 ( .gnd(gnd), .vdd(vdd), .A(_2529_), .B(_2530_), .C(_2531_), .Y(_2533_) );
NAND3X1 NAND3X1_423 ( .gnd(gnd), .vdd(vdd), .A(_2528_), .B(_2533_), .C(_2270_), .Y(_2534_) );
AOI21X1 AOI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_2166_), .B(_1911_), .C(_2171_), .Y(_2535_) );
AOI21X1 AOI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_2530_), .B(_2531_), .C(_2529_), .Y(_2536_) );
AOI21X1 AOI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .B(_2527_), .C(_2157_), .Y(_2537_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_2536_), .B(_2537_), .C(_2535_), .Y(_2538_) );
NAND3X1 NAND3X1_424 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .B(_2538_), .C(_2534_), .Y(_2539_) );
NOR3X1 NOR3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_2536_), .B(_2535_), .C(_2537_), .Y(_2540_) );
AOI21X1 AOI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_2528_), .B(_2533_), .C(_2270_), .Y(_2541_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_2540_), .B(_2541_), .C(_3224_), .Y(_2542_) );
NAND3X1 NAND3X1_425 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_2539_), .C(_2542_), .Y(_2544_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_2269_), .B(_2544_), .Y(_2545_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_2540_), .B(_2541_), .C(_3222_), .Y(_2546_) );
NAND3X1 NAND3X1_426 ( .gnd(gnd), .vdd(vdd), .A(_3224_), .B(_2538_), .C(_2534_), .Y(_2547_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .B(_2546_), .Y(_2548_) );
NAND3X1 NAND3X1_427 ( .gnd(gnd), .vdd(vdd), .A(W_205_), .B(_394_), .C(_2548_), .Y(_2549_) );
AOI21X1 AOI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .B(_2549_), .C(_2267_), .Y(_2550_) );
NAND3X1 NAND3X1_428 ( .gnd(gnd), .vdd(vdd), .A(_2269_), .B(_394_), .C(_2548_), .Y(_2551_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(W_205_), .B(_2544_), .Y(_2552_) );
AOI21X1 AOI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2552_), .C(_2179_), .Y(_2553_) );
NOR3X1 NOR3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_2550_), .B(_2266_), .C(_2553_), .Y(_2555_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_2191_), .B(_2194_), .C(_2185_), .Y(_2556_) );
NAND3X1 NAND3X1_429 ( .gnd(gnd), .vdd(vdd), .A(_2179_), .B(_2551_), .C(_2552_), .Y(_2557_) );
NAND3X1 NAND3X1_430 ( .gnd(gnd), .vdd(vdd), .A(_2267_), .B(_2545_), .C(_2549_), .Y(_2558_) );
AOI21X1 AOI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_2557_), .B(_2558_), .C(_2556_), .Y(_2559_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_2555_), .B(_2559_), .C(_3230_), .Y(_2560_) );
NAND3X1 NAND3X1_431 ( .gnd(gnd), .vdd(vdd), .A(_2557_), .B(_2558_), .C(_2556_), .Y(_2561_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_2550_), .B(_2553_), .C(_2266_), .Y(_2562_) );
NAND3X1 NAND3X1_432 ( .gnd(gnd), .vdd(vdd), .A(_3232_), .B(_2562_), .C(_2561_), .Y(_2563_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_2563_), .B(_2560_), .Y(_2564_) );
NAND3X1 NAND3X1_433 ( .gnd(gnd), .vdd(vdd), .A(_2265_), .B(_402_), .C(_2564_), .Y(_2566_) );
NAND3X1 NAND3X1_434 ( .gnd(gnd), .vdd(vdd), .A(_3230_), .B(_2562_), .C(_2561_), .Y(_2567_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_2555_), .B(_2559_), .C(_3232_), .Y(_2568_) );
NAND3X1 NAND3X1_435 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_2567_), .C(_2568_), .Y(_2569_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(W_221_), .B(_2569_), .Y(_2570_) );
NAND3X1 NAND3X1_436 ( .gnd(gnd), .vdd(vdd), .A(_2204_), .B(_2566_), .C(_2570_), .Y(_2571_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(_2204_), .Y(_2572_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_2265_), .B(_2569_), .Y(_2573_) );
NAND3X1 NAND3X1_437 ( .gnd(gnd), .vdd(vdd), .A(W_221_), .B(_402_), .C(_2564_), .Y(_2574_) );
NAND3X1 NAND3X1_438 ( .gnd(gnd), .vdd(vdd), .A(_2572_), .B(_2573_), .C(_2574_), .Y(_2575_) );
NAND3X1 NAND3X1_439 ( .gnd(gnd), .vdd(vdd), .A(_2571_), .B(_2575_), .C(_2264_), .Y(_2577_) );
AOI21X1 AOI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_2211_), .B(_1908_), .C(_2215_), .Y(_2578_) );
AOI21X1 AOI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_2573_), .B(_2574_), .C(_2572_), .Y(_2579_) );
AOI21X1 AOI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_2566_), .B(_2570_), .C(_2204_), .Y(_2580_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_2579_), .B(_2580_), .C(_2578_), .Y(_2581_) );
AOI21X1 AOI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_2577_), .B(_2581_), .C(_3238_), .Y(_2582_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(_2582_), .Y(_2583_) );
NAND3X1 NAND3X1_440 ( .gnd(gnd), .vdd(vdd), .A(_3238_), .B(_2577_), .C(_2581_), .Y(_2584_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_2584_), .B(_410_), .Y(_2585_) );
NAND3X1 NAND3X1_441 ( .gnd(gnd), .vdd(vdd), .A(_2263_), .B(_2583_), .C(_2585_), .Y(_2586_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_2584_), .Y(_2588_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .B(_2582_), .C(W_237_), .Y(_2589_) );
NAND3X1 NAND3X1_442 ( .gnd(gnd), .vdd(vdd), .A(_2226_), .B(_2589_), .C(_2586_), .Y(_2590_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(_2226_), .Y(_2591_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .B(_2582_), .C(_2263_), .Y(_2592_) );
NAND3X1 NAND3X1_443 ( .gnd(gnd), .vdd(vdd), .A(W_237_), .B(_2583_), .C(_2585_), .Y(_2593_) );
NAND3X1 NAND3X1_444 ( .gnd(gnd), .vdd(vdd), .A(_2591_), .B(_2592_), .C(_2593_), .Y(_2594_) );
NAND3X1 NAND3X1_445 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .B(_2594_), .C(_2262_), .Y(_2595_) );
AOI21X1 AOI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_2235_), .B(_1905_), .C(_2239_), .Y(_2596_) );
AOI21X1 AOI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_2592_), .B(_2593_), .C(_2591_), .Y(_2597_) );
AOI21X1 AOI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_2589_), .B(_2586_), .C(_2226_), .Y(_2599_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_2597_), .B(_2599_), .C(_2596_), .Y(_2600_) );
NAND3X1 NAND3X1_446 ( .gnd(gnd), .vdd(vdd), .A(_3247_), .B(_2595_), .C(_2600_), .Y(_2601_) );
NOR3X1 NOR3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_2597_), .B(_2599_), .C(_2596_), .Y(_2602_) );
AOI21X1 AOI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .B(_2594_), .C(_2262_), .Y(_2603_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_2602_), .B(_2603_), .C(_3249_), .Y(_2604_) );
NAND3X1 NAND3X1_447 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_2601_), .C(_2604_), .Y(_2605_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_2261_), .B(_2605_), .Y(_2606_) );
NAND3X1 NAND3X1_448 ( .gnd(gnd), .vdd(vdd), .A(_3249_), .B(_2595_), .C(_2600_), .Y(_2607_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2602_), .B(_2603_), .C(_3247_), .Y(_2608_) );
AOI21X1 AOI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_2607_), .B(_2608_), .C(_418_), .Y(_2610_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(W_253_), .B(_2610_), .Y(_2611_) );
AOI21X1 AOI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_2606_), .B(_2611_), .C(_2260_), .Y(_2612_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(_2612_), .Y(_2613_) );
NAND3X1 NAND3X1_449 ( .gnd(gnd), .vdd(vdd), .A(_2260_), .B(_2606_), .C(_2611_), .Y(_2614_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_2614_), .B(_2613_), .Y(_2615_) );
XNOR2X1 XNOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_2615_), .B(_2258_), .Y(H_21_) );
AOI21X1 AOI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_2258_), .B(_2614_), .C(_2612_), .Y(_2616_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(W_253_), .B(_2605_), .Y(_2617_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(W_254_), .Y(_2618_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_2596_), .B(_2597_), .C(_2594_), .Y(_2620_) );
AOI21X1 AOI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_2571_), .B(_2264_), .C(_2580_), .Y(_2621_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(_2566_), .Y(_2622_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(W_222_), .Y(_2623_) );
AOI21X1 AOI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_2557_), .B(_2556_), .C(_2553_), .Y(_2624_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .Y(_2625_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(W_206_), .Y(_2626_) );
AOI21X1 AOI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_2528_), .B(_2270_), .C(_2537_), .Y(_2627_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(W_190_), .Y(_2628_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2514_), .B(_2513_), .C(_2511_), .Y(_2629_) );
AOI21X1 AOI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_2275_), .B(_2484_), .C(_2493_), .Y(_2631_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(_2631_), .Y(_2632_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .B(_2469_), .C(_2467_), .Y(_2633_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_2449_), .B(_2443_), .Y(_2634_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[94]), .Y(_2635_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_2426_), .B(_2420_), .Y(_2636_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_2403_), .B(_2397_), .Y(_2637_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_2379_), .B(_2373_), .Y(_2638_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_2358_), .B(_2363_), .Y(_2639_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(_2639_), .Y(_2640_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_2328_), .B(_2333_), .Y(_2642_) );
INVX2 INVX2_45 ( .gnd(gnd), .vdd(vdd), .A(_2642_), .Y(_2643_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[14]), .Y(_2644_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_2289_), .B(_2307_), .C(_2313_), .Y(_2645_) );
INVX2 INVX2_46 ( .gnd(gnd), .vdd(vdd), .A(_2645_), .Y(_2646_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(W_30_), .Y(_2647_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(W_12_), .B(W_13_), .Y(_2648_) );
XNOR2X1 XNOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_2648_), .B(W_14_), .Y(_2649_) );
XNOR2X1 XNOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_809_), .B(W_10_), .Y(_2650_) );
XNOR2X1 XNOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_2650_), .B(_2649_), .Y(_2651_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_2651_), .B(_2647_), .Y(_2653_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_2647_), .B(_2651_), .Y(_2654_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_2654_), .B(_2653_), .Y(_2655_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_2655_), .B(_2305_), .Y(_2656_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_2305_), .B(_2655_), .Y(_2657_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_2657_), .B(_2656_), .Y(_2658_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_2646_), .B(_2658_), .Y(_2659_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_2656_), .B(_2657_), .Y(_2660_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_2304_), .B(_2320_), .C(_2660_), .Y(_2661_) );
XNOR2X1 XNOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_823_), .B(_855_), .Y(_2662_) );
NAND3X1 NAND3X1_450 ( .gnd(gnd), .vdd(vdd), .A(_2659_), .B(_2662_), .C(_2661_), .Y(_2664_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_2645_), .B(_2660_), .Y(_2665_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_2646_), .B(_2658_), .Y(_2666_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(_2662_), .Y(_2667_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_2665_), .B(_2666_), .C(_2667_), .Y(_2668_) );
NAND3X1 NAND3X1_451 ( .gnd(gnd), .vdd(vdd), .A(_2644_), .B(_2664_), .C(_2668_), .Y(_2669_) );
NAND3X1 NAND3X1_452 ( .gnd(gnd), .vdd(vdd), .A(_2659_), .B(_2667_), .C(_2661_), .Y(_2670_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_2665_), .B(_2666_), .C(_2662_), .Y(_2671_) );
NAND3X1 NAND3X1_453 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[14]), .B(_2670_), .C(_2671_), .Y(_2672_) );
AOI21X1 AOI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_2669_), .B(_2672_), .C(_2322_), .Y(_2673_) );
NAND3X1 NAND3X1_454 ( .gnd(gnd), .vdd(vdd), .A(_2322_), .B(_2669_), .C(_2672_), .Y(_2675_) );
INVX2 INVX2_47 ( .gnd(gnd), .vdd(vdd), .A(_2675_), .Y(_2676_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_2676_), .B(_2673_), .C(_2643_), .Y(_2677_) );
INVX2 INVX2_48 ( .gnd(gnd), .vdd(vdd), .A(_2673_), .Y(_2678_) );
NAND3X1 NAND3X1_455 ( .gnd(gnd), .vdd(vdd), .A(_2642_), .B(_2675_), .C(_2678_), .Y(_2679_) );
XNOR2X1 XNOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_887_), .B(_844_), .Y(_2680_) );
NAND3X1 NAND3X1_456 ( .gnd(gnd), .vdd(vdd), .A(_2680_), .B(_2679_), .C(_2677_), .Y(_2681_) );
AOI21X1 AOI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_2675_), .B(_2678_), .C(_2642_), .Y(_2682_) );
NOR3X1 NOR3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_2673_), .B(_2643_), .C(_2676_), .Y(_2683_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(_2680_), .Y(_2684_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2682_), .C(_2684_), .Y(_2686_) );
NAND3X1 NAND3X1_457 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[30]), .B(_2681_), .C(_2686_), .Y(_2687_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[30]), .Y(_2688_) );
NAND3X1 NAND3X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2684_), .B(_2679_), .C(_2677_), .Y(_2689_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2682_), .C(_2680_), .Y(_2690_) );
NAND3X1 NAND3X1_459 ( .gnd(gnd), .vdd(vdd), .A(_2688_), .B(_2689_), .C(_2690_), .Y(_2691_) );
NAND3X1 NAND3X1_460 ( .gnd(gnd), .vdd(vdd), .A(_2352_), .B(_2687_), .C(_2691_), .Y(_2692_) );
NAND3X1 NAND3X1_461 ( .gnd(gnd), .vdd(vdd), .A(_2688_), .B(_2681_), .C(_2686_), .Y(_2693_) );
NAND3X1 NAND3X1_462 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[30]), .B(_2689_), .C(_2690_), .Y(_2694_) );
NAND3X1 NAND3X1_463 ( .gnd(gnd), .vdd(vdd), .A(_2346_), .B(_2693_), .C(_2694_), .Y(_2695_) );
NAND3X1 NAND3X1_464 ( .gnd(gnd), .vdd(vdd), .A(_2640_), .B(_2692_), .C(_2695_), .Y(_2697_) );
NAND3X1 NAND3X1_465 ( .gnd(gnd), .vdd(vdd), .A(_2346_), .B(_2687_), .C(_2691_), .Y(_2698_) );
NAND3X1 NAND3X1_466 ( .gnd(gnd), .vdd(vdd), .A(_2352_), .B(_2693_), .C(_2694_), .Y(_2699_) );
NAND3X1 NAND3X1_467 ( .gnd(gnd), .vdd(vdd), .A(_2639_), .B(_2698_), .C(_2699_), .Y(_2700_) );
XNOR2X1 XNOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_925_), .B(_876_), .Y(_2701_) );
NAND3X1 NAND3X1_468 ( .gnd(gnd), .vdd(vdd), .A(_2701_), .B(_2697_), .C(_2700_), .Y(_2702_) );
AOI21X1 AOI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_2698_), .B(_2699_), .C(_2639_), .Y(_2703_) );
AOI21X1 AOI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_2692_), .B(_2695_), .C(_2640_), .Y(_2704_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(_2701_), .Y(_2705_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_2703_), .B(_2704_), .C(_2705_), .Y(_2706_) );
NAND3X1 NAND3X1_469 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[46]), .B(_2702_), .C(_2706_), .Y(_2708_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[46]), .Y(_2709_) );
NAND3X1 NAND3X1_470 ( .gnd(gnd), .vdd(vdd), .A(_2705_), .B(_2697_), .C(_2700_), .Y(_2710_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_2703_), .B(_2704_), .C(_2701_), .Y(_2711_) );
NAND3X1 NAND3X1_471 ( .gnd(gnd), .vdd(vdd), .A(_2709_), .B(_2710_), .C(_2711_), .Y(_2712_) );
NAND3X1 NAND3X1_472 ( .gnd(gnd), .vdd(vdd), .A(_2368_), .B(_2708_), .C(_2712_), .Y(_2713_) );
NAND3X1 NAND3X1_473 ( .gnd(gnd), .vdd(vdd), .A(_2709_), .B(_2702_), .C(_2706_), .Y(_2714_) );
NAND3X1 NAND3X1_474 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[46]), .B(_2710_), .C(_2711_), .Y(_2715_) );
NAND3X1 NAND3X1_475 ( .gnd(gnd), .vdd(vdd), .A(_2375_), .B(_2714_), .C(_2715_), .Y(_2716_) );
NAND3X1 NAND3X1_476 ( .gnd(gnd), .vdd(vdd), .A(_2638_), .B(_2713_), .C(_2716_), .Y(_2717_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_2373_), .B(_2379_), .Y(_2719_) );
NAND3X1 NAND3X1_477 ( .gnd(gnd), .vdd(vdd), .A(_2375_), .B(_2708_), .C(_2712_), .Y(_2720_) );
NAND3X1 NAND3X1_478 ( .gnd(gnd), .vdd(vdd), .A(_2368_), .B(_2714_), .C(_2715_), .Y(_2721_) );
NAND3X1 NAND3X1_479 ( .gnd(gnd), .vdd(vdd), .A(_2719_), .B(_2720_), .C(_2721_), .Y(_2722_) );
XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_960_), .B(_910_), .Y(_2723_) );
NAND3X1 NAND3X1_480 ( .gnd(gnd), .vdd(vdd), .A(_2723_), .B(_2722_), .C(_2717_), .Y(_2724_) );
AOI21X1 AOI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_2720_), .B(_2721_), .C(_2719_), .Y(_2725_) );
AOI21X1 AOI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_2713_), .B(_2716_), .C(_2638_), .Y(_2726_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(_2723_), .Y(_2727_) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_2726_), .B(_2725_), .C(_2727_), .Y(_2728_) );
NAND3X1 NAND3X1_481 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[62]), .B(_2724_), .C(_2728_), .Y(_2730_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[62]), .Y(_2731_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2726_), .B(_2725_), .C(_2723_), .Y(_2732_) );
NAND3X1 NAND3X1_482 ( .gnd(gnd), .vdd(vdd), .A(_2727_), .B(_2722_), .C(_2717_), .Y(_2733_) );
NAND3X1 NAND3X1_483 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .B(_2733_), .C(_2732_), .Y(_2734_) );
NAND3X1 NAND3X1_484 ( .gnd(gnd), .vdd(vdd), .A(_2392_), .B(_2730_), .C(_2734_), .Y(_2735_) );
NAND3X1 NAND3X1_485 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .B(_2724_), .C(_2728_), .Y(_2736_) );
NAND3X1 NAND3X1_486 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[62]), .B(_2733_), .C(_2732_), .Y(_2737_) );
NAND3X1 NAND3X1_487 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .B(_2736_), .C(_2737_), .Y(_2738_) );
NAND3X1 NAND3X1_488 ( .gnd(gnd), .vdd(vdd), .A(_2735_), .B(_2738_), .C(_2637_), .Y(_2739_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_2397_), .B(_2403_), .Y(_2741_) );
NAND3X1 NAND3X1_489 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .B(_2730_), .C(_2734_), .Y(_2742_) );
NAND3X1 NAND3X1_490 ( .gnd(gnd), .vdd(vdd), .A(_2392_), .B(_2736_), .C(_2737_), .Y(_2743_) );
NAND3X1 NAND3X1_491 ( .gnd(gnd), .vdd(vdd), .A(_2741_), .B(_2742_), .C(_2743_), .Y(_2744_) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_3346_), .B(_3349_), .C(_1001_), .Y(_2745_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .B(_997_), .C(_962_), .Y(_2746_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_2746_), .B(_2745_), .Y(_2747_) );
NAND3X1 NAND3X1_492 ( .gnd(gnd), .vdd(vdd), .A(_2747_), .B(_2744_), .C(_2739_), .Y(_2748_) );
AOI21X1 AOI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_2742_), .B(_2743_), .C(_2741_), .Y(_2749_) );
AOI21X1 AOI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_2735_), .B(_2738_), .C(_2637_), .Y(_2750_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(_2747_), .Y(_2752_) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_2750_), .B(_2749_), .C(_2752_), .Y(_2753_) );
NAND3X1 NAND3X1_493 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[78]), .B(_2748_), .C(_2753_), .Y(_2754_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[78]), .Y(_2755_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_2750_), .B(_2749_), .C(_2747_), .Y(_2756_) );
NAND3X1 NAND3X1_494 ( .gnd(gnd), .vdd(vdd), .A(_2752_), .B(_2744_), .C(_2739_), .Y(_2757_) );
NAND3X1 NAND3X1_495 ( .gnd(gnd), .vdd(vdd), .A(_2755_), .B(_2757_), .C(_2756_), .Y(_2758_) );
NAND3X1 NAND3X1_496 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .B(_2754_), .C(_2758_), .Y(_2759_) );
NAND3X1 NAND3X1_497 ( .gnd(gnd), .vdd(vdd), .A(_2755_), .B(_2748_), .C(_2753_), .Y(_2760_) );
NAND3X1 NAND3X1_498 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[78]), .B(_2757_), .C(_2756_), .Y(_2761_) );
NAND3X1 NAND3X1_499 ( .gnd(gnd), .vdd(vdd), .A(_2423_), .B(_2760_), .C(_2761_), .Y(_2763_) );
NAND3X1 NAND3X1_500 ( .gnd(gnd), .vdd(vdd), .A(_2759_), .B(_2763_), .C(_2636_), .Y(_2764_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_2420_), .B(_2426_), .Y(_2765_) );
NAND3X1 NAND3X1_501 ( .gnd(gnd), .vdd(vdd), .A(_2423_), .B(_2754_), .C(_2758_), .Y(_2766_) );
NAND3X1 NAND3X1_502 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .B(_2760_), .C(_2761_), .Y(_2767_) );
NAND3X1 NAND3X1_503 ( .gnd(gnd), .vdd(vdd), .A(_2766_), .B(_2767_), .C(_2765_), .Y(_2768_) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_3358_), .B(_3361_), .C(_1045_), .Y(_2769_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(_2769_), .Y(_2770_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .Y(_2771_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_2771_), .B(_1045_), .Y(_2772_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_2772_), .B(_2770_), .Y(_2774_) );
NAND3X1 NAND3X1_504 ( .gnd(gnd), .vdd(vdd), .A(_2774_), .B(_2768_), .C(_2764_), .Y(_2775_) );
AOI21X1 AOI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_2766_), .B(_2767_), .C(_2765_), .Y(_2776_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_2420_), .B(_2426_), .C(_2759_), .D(_2763_), .Y(_2777_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(_2774_), .Y(_2778_) );
OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_2777_), .B(_2776_), .C(_2778_), .Y(_2779_) );
NAND3X1 NAND3X1_505 ( .gnd(gnd), .vdd(vdd), .A(_2635_), .B(_2779_), .C(_2775_), .Y(_2780_) );
NAND3X1 NAND3X1_506 ( .gnd(gnd), .vdd(vdd), .A(_2778_), .B(_2768_), .C(_2764_), .Y(_2781_) );
OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_2777_), .B(_2776_), .C(_2774_), .Y(_2782_) );
NAND3X1 NAND3X1_507 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[94]), .B(_2782_), .C(_2781_), .Y(_2783_) );
AOI21X1 AOI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_2780_), .B(_2783_), .C(_2438_), .Y(_2785_) );
NAND3X1 NAND3X1_508 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[94]), .B(_2779_), .C(_2775_), .Y(_2786_) );
NAND3X1 NAND3X1_509 ( .gnd(gnd), .vdd(vdd), .A(_2635_), .B(_2782_), .C(_2781_), .Y(_2787_) );
AOI21X1 AOI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_2786_), .B(_2787_), .C(_2446_), .Y(_2788_) );
OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_2785_), .B(_2788_), .C(_2634_), .Y(_2789_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_2443_), .B(_2449_), .Y(_2790_) );
NAND3X1 NAND3X1_510 ( .gnd(gnd), .vdd(vdd), .A(_2446_), .B(_2786_), .C(_2787_), .Y(_2791_) );
NAND3X1 NAND3X1_511 ( .gnd(gnd), .vdd(vdd), .A(_2438_), .B(_2780_), .C(_2783_), .Y(_2792_) );
NAND3X1 NAND3X1_512 ( .gnd(gnd), .vdd(vdd), .A(_2791_), .B(_2792_), .C(_2790_), .Y(_2793_) );
AOI21X1 AOI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_2793_), .B(_2789_), .C(_1028_), .Y(_2794_) );
NAND3X1 NAND3X1_513 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_2793_), .C(_2789_), .Y(_2796_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1075_), .B(_2796_), .Y(_2797_) );
OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_2797_), .B(_2794_), .C(W_142_), .Y(_2798_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(W_142_), .Y(_2799_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(_2794_), .Y(_2800_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_2796_), .B(_1075_), .Y(_2801_) );
NAND3X1 NAND3X1_514 ( .gnd(gnd), .vdd(vdd), .A(_2799_), .B(_2800_), .C(_2801_), .Y(_2802_) );
NAND3X1 NAND3X1_515 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .B(_2798_), .C(_2802_), .Y(_2803_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .Y(_2804_) );
OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_2797_), .B(_2794_), .C(_2799_), .Y(_2805_) );
NAND3X1 NAND3X1_516 ( .gnd(gnd), .vdd(vdd), .A(W_142_), .B(_2800_), .C(_2801_), .Y(_2807_) );
NAND3X1 NAND3X1_517 ( .gnd(gnd), .vdd(vdd), .A(_2804_), .B(_2805_), .C(_2807_), .Y(_2808_) );
AOI21X1 AOI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_2803_), .B(_2808_), .C(_2633_), .Y(_2809_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(_2633_), .Y(_2810_) );
NAND3X1 NAND3X1_518 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .B(_2805_), .C(_2807_), .Y(_2811_) );
NAND3X1 NAND3X1_519 ( .gnd(gnd), .vdd(vdd), .A(_2804_), .B(_2798_), .C(_2802_), .Y(_2812_) );
AOI21X1 AOI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_2811_), .B(_2812_), .C(_2810_), .Y(_2813_) );
OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_2809_), .B(_2813_), .C(_789_), .Y(_2814_) );
NAND3X1 NAND3X1_520 ( .gnd(gnd), .vdd(vdd), .A(_2810_), .B(_2811_), .C(_2812_), .Y(_2815_) );
NAND3X1 NAND3X1_521 ( .gnd(gnd), .vdd(vdd), .A(_2633_), .B(_2803_), .C(_2808_), .Y(_2816_) );
NAND3X1 NAND3X1_522 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_2816_), .C(_2815_), .Y(_2818_) );
NAND3X1 NAND3X1_523 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(_2818_), .C(_2814_), .Y(_2819_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(W_158_), .B(_2819_), .Y(_2820_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(W_158_), .Y(_2821_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_2818_), .B(_1105_), .Y(_2822_) );
NAND3X1 NAND3X1_524 ( .gnd(gnd), .vdd(vdd), .A(_2821_), .B(_2814_), .C(_2822_), .Y(_2823_) );
NAND3X1 NAND3X1_525 ( .gnd(gnd), .vdd(vdd), .A(_2479_), .B(_2820_), .C(_2823_), .Y(_2824_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(_2479_), .Y(_2825_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_2821_), .B(_2819_), .Y(_2826_) );
NAND3X1 NAND3X1_526 ( .gnd(gnd), .vdd(vdd), .A(W_158_), .B(_2814_), .C(_2822_), .Y(_2827_) );
NAND3X1 NAND3X1_527 ( .gnd(gnd), .vdd(vdd), .A(_2825_), .B(_2826_), .C(_2827_), .Y(_2829_) );
AOI21X1 AOI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_2824_), .B(_2829_), .C(_2632_), .Y(_2830_) );
NAND3X1 NAND3X1_528 ( .gnd(gnd), .vdd(vdd), .A(_2479_), .B(_2826_), .C(_2827_), .Y(_2831_) );
NAND3X1 NAND3X1_529 ( .gnd(gnd), .vdd(vdd), .A(_2825_), .B(_2820_), .C(_2823_), .Y(_2832_) );
AOI21X1 AOI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_2831_), .B(_2832_), .C(_2631_), .Y(_2833_) );
OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_2830_), .B(_2833_), .C(_784_), .Y(_2834_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(_2834_), .Y(_2835_) );
NAND3X1 NAND3X1_530 ( .gnd(gnd), .vdd(vdd), .A(_2631_), .B(_2831_), .C(_2832_), .Y(_2836_) );
NAND3X1 NAND3X1_531 ( .gnd(gnd), .vdd(vdd), .A(_2824_), .B(_2632_), .C(_2829_), .Y(_2837_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_2836_), .B(_2837_), .Y(_2838_) );
OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2838_), .B(_784_), .C(_1136_), .Y(_2840_) );
OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_2840_), .B(_2835_), .C(W_174_), .Y(_2841_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(W_174_), .Y(_2842_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_2830_), .B(_2833_), .Y(_2843_) );
AOI21X1 AOI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_2843_), .C(_1140_), .Y(_2844_) );
NAND3X1 NAND3X1_532 ( .gnd(gnd), .vdd(vdd), .A(_2842_), .B(_2834_), .C(_2844_), .Y(_2845_) );
NAND3X1 NAND3X1_533 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .B(_2841_), .C(_2845_), .Y(_2846_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .Y(_2847_) );
OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_2840_), .B(_2835_), .C(_2842_), .Y(_2848_) );
NAND3X1 NAND3X1_534 ( .gnd(gnd), .vdd(vdd), .A(W_174_), .B(_2834_), .C(_2844_), .Y(_2849_) );
NAND3X1 NAND3X1_535 ( .gnd(gnd), .vdd(vdd), .A(_2847_), .B(_2848_), .C(_2849_), .Y(_2851_) );
AOI21X1 AOI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_2846_), .B(_2851_), .C(_2629_), .Y(_2852_) );
AOI21X1 AOI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_2272_), .B(_2506_), .C(_2515_), .Y(_2853_) );
NAND3X1 NAND3X1_536 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .B(_2848_), .C(_2849_), .Y(_2854_) );
NAND3X1 NAND3X1_537 ( .gnd(gnd), .vdd(vdd), .A(_2847_), .B(_2841_), .C(_2845_), .Y(_2855_) );
AOI21X1 AOI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_2854_), .B(_2855_), .C(_2853_), .Y(_2856_) );
OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_2852_), .B(_2856_), .C(_779_), .Y(_2857_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .Y(_2858_) );
NAND3X1 NAND3X1_538 ( .gnd(gnd), .vdd(vdd), .A(_2853_), .B(_2854_), .C(_2855_), .Y(_2859_) );
NAND3X1 NAND3X1_539 ( .gnd(gnd), .vdd(vdd), .A(_2629_), .B(_2846_), .C(_2851_), .Y(_2860_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_2859_), .B(_2860_), .Y(_2862_) );
OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_2862_), .B(_779_), .C(_1169_), .Y(_2863_) );
OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_2863_), .B(_2858_), .C(_2628_), .Y(_2864_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_2852_), .B(_2856_), .Y(_2865_) );
AOI21X1 AOI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_2865_), .C(_1173_), .Y(_2866_) );
NAND3X1 NAND3X1_540 ( .gnd(gnd), .vdd(vdd), .A(W_190_), .B(_2857_), .C(_2866_), .Y(_2867_) );
NAND3X1 NAND3X1_541 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .B(_2864_), .C(_2867_), .Y(_2868_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .Y(_2869_) );
OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_2863_), .B(_2858_), .C(W_190_), .Y(_2870_) );
NAND3X1 NAND3X1_542 ( .gnd(gnd), .vdd(vdd), .A(_2628_), .B(_2857_), .C(_2866_), .Y(_2871_) );
NAND3X1 NAND3X1_543 ( .gnd(gnd), .vdd(vdd), .A(_2869_), .B(_2870_), .C(_2871_), .Y(_2873_) );
NAND3X1 NAND3X1_544 ( .gnd(gnd), .vdd(vdd), .A(_2627_), .B(_2868_), .C(_2873_), .Y(_2874_) );
OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_2536_), .B(_2535_), .C(_2533_), .Y(_2875_) );
NAND3X1 NAND3X1_545 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .B(_2870_), .C(_2871_), .Y(_2876_) );
NAND3X1 NAND3X1_546 ( .gnd(gnd), .vdd(vdd), .A(_2869_), .B(_2864_), .C(_2867_), .Y(_2877_) );
NAND3X1 NAND3X1_547 ( .gnd(gnd), .vdd(vdd), .A(_2875_), .B(_2876_), .C(_2877_), .Y(_2878_) );
NAND3X1 NAND3X1_548 ( .gnd(gnd), .vdd(vdd), .A(_775_), .B(_2878_), .C(_2874_), .Y(_2879_) );
AOI21X1 AOI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_2876_), .B(_2877_), .C(_2875_), .Y(_2880_) );
AOI21X1 AOI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_2868_), .B(_2873_), .C(_2627_), .Y(_2881_) );
OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_2880_), .B(_2881_), .C(_774_), .Y(_2882_) );
NAND3X1 NAND3X1_549 ( .gnd(gnd), .vdd(vdd), .A(_1202_), .B(_2879_), .C(_2882_), .Y(_2884_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_2626_), .B(_2884_), .Y(_2885_) );
OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_2880_), .B(_2881_), .C(_775_), .Y(_2886_) );
NAND3X1 NAND3X1_550 ( .gnd(gnd), .vdd(vdd), .A(_774_), .B(_2878_), .C(_2874_), .Y(_2887_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_2887_), .B(_2886_), .Y(_2888_) );
NAND3X1 NAND3X1_551 ( .gnd(gnd), .vdd(vdd), .A(W_206_), .B(_1202_), .C(_2888_), .Y(_2889_) );
AOI21X1 AOI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_2889_), .B(_2885_), .C(_2625_), .Y(_2890_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(W_206_), .B(_2884_), .Y(_2891_) );
NAND3X1 NAND3X1_552 ( .gnd(gnd), .vdd(vdd), .A(_2626_), .B(_1202_), .C(_2888_), .Y(_2892_) );
AOI21X1 AOI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_2892_), .B(_2891_), .C(_2551_), .Y(_2893_) );
OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2890_), .B(_2893_), .C(_2624_), .Y(_2895_) );
OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2550_), .B(_2266_), .C(_2558_), .Y(_2896_) );
NAND3X1 NAND3X1_553 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2892_), .C(_2891_), .Y(_2897_) );
NAND3X1 NAND3X1_554 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .B(_2889_), .C(_2885_), .Y(_2898_) );
NAND3X1 NAND3X1_555 ( .gnd(gnd), .vdd(vdd), .A(_2896_), .B(_2897_), .C(_2898_), .Y(_2899_) );
AOI21X1 AOI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_2899_), .B(_2895_), .C(_1209_), .Y(_2900_) );
NAND3X1 NAND3X1_556 ( .gnd(gnd), .vdd(vdd), .A(_1209_), .B(_2899_), .C(_2895_), .Y(_2901_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1234_), .B(_2901_), .Y(_2902_) );
OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2902_), .B(_2900_), .C(_2623_), .Y(_2903_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(_2900_), .Y(_2904_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_2901_), .B(_1234_), .Y(_2906_) );
NAND3X1 NAND3X1_557 ( .gnd(gnd), .vdd(vdd), .A(W_222_), .B(_2904_), .C(_2906_), .Y(_2907_) );
AOI21X1 AOI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_2903_), .B(_2907_), .C(_2622_), .Y(_2908_) );
OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_2902_), .B(_2900_), .C(W_222_), .Y(_2909_) );
NAND3X1 NAND3X1_558 ( .gnd(gnd), .vdd(vdd), .A(_2623_), .B(_2904_), .C(_2906_), .Y(_2910_) );
AOI21X1 AOI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_2909_), .B(_2910_), .C(_2566_), .Y(_2911_) );
OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_2908_), .B(_2911_), .C(_2621_), .Y(_2912_) );
OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_2578_), .B(_2579_), .C(_2575_), .Y(_2913_) );
NAND3X1 NAND3X1_559 ( .gnd(gnd), .vdd(vdd), .A(_2566_), .B(_2909_), .C(_2910_), .Y(_2914_) );
NAND3X1 NAND3X1_560 ( .gnd(gnd), .vdd(vdd), .A(_2622_), .B(_2903_), .C(_2907_), .Y(_2915_) );
NAND3X1 NAND3X1_561 ( .gnd(gnd), .vdd(vdd), .A(_2914_), .B(_2915_), .C(_2913_), .Y(_2917_) );
AOI21X1 AOI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_2917_), .B(_2912_), .C(_767_), .Y(_2918_) );
NAND3X1 NAND3X1_562 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_2917_), .C(_2912_), .Y(_2919_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1270_), .B(_2919_), .Y(_2920_) );
OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_2920_), .B(_2918_), .C(W_238_), .Y(_2921_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(W_238_), .Y(_2922_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(_2918_), .Y(_2923_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_2919_), .B(_1270_), .Y(_2924_) );
NAND3X1 NAND3X1_563 ( .gnd(gnd), .vdd(vdd), .A(_2922_), .B(_2923_), .C(_2924_), .Y(_2925_) );
NAND3X1 NAND3X1_564 ( .gnd(gnd), .vdd(vdd), .A(_2586_), .B(_2921_), .C(_2925_), .Y(_2926_) );
INVX2 INVX2_49 ( .gnd(gnd), .vdd(vdd), .A(_2586_), .Y(_2928_) );
OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_2920_), .B(_2918_), .C(_2922_), .Y(_2929_) );
NAND3X1 NAND3X1_565 ( .gnd(gnd), .vdd(vdd), .A(W_238_), .B(_2923_), .C(_2924_), .Y(_2930_) );
NAND3X1 NAND3X1_566 ( .gnd(gnd), .vdd(vdd), .A(_2928_), .B(_2929_), .C(_2930_), .Y(_2931_) );
AOI21X1 AOI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .B(_2931_), .C(_2620_), .Y(_2932_) );
AOI21X1 AOI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .B(_2262_), .C(_2599_), .Y(_2933_) );
NAND3X1 NAND3X1_567 ( .gnd(gnd), .vdd(vdd), .A(_2586_), .B(_2929_), .C(_2930_), .Y(_2934_) );
NAND3X1 NAND3X1_568 ( .gnd(gnd), .vdd(vdd), .A(_2928_), .B(_2921_), .C(_2925_), .Y(_2935_) );
AOI21X1 AOI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_2934_), .B(_2935_), .C(_2933_), .Y(_2936_) );
OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_2932_), .B(_2936_), .C(_3456_), .Y(_2937_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(_2937_), .Y(_2939_) );
AOI21X1 AOI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_2929_), .B(_2930_), .C(_2928_), .Y(_2940_) );
AOI21X1 AOI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_2921_), .B(_2925_), .C(_2586_), .Y(_2941_) );
OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_2940_), .B(_2941_), .C(_2933_), .Y(_2942_) );
NAND3X1 NAND3X1_569 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .B(_2931_), .C(_2620_), .Y(_2943_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_2943_), .B(_2942_), .Y(_2944_) );
OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_2944_), .B(_3456_), .C(_1306_), .Y(_2945_) );
OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_2945_), .B(_2939_), .C(_2618_), .Y(_2946_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_2932_), .B(_2936_), .Y(_2947_) );
AOI21X1 AOI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_3457_), .B(_2947_), .C(_1307_), .Y(_2948_) );
NAND3X1 NAND3X1_570 ( .gnd(gnd), .vdd(vdd), .A(W_254_), .B(_2937_), .C(_2948_), .Y(_2950_) );
AOI21X1 AOI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2950_), .B(_2946_), .C(_2617_), .Y(_2951_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(_2617_), .Y(_2952_) );
OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_2945_), .B(_2939_), .C(W_254_), .Y(_2953_) );
NAND3X1 NAND3X1_571 ( .gnd(gnd), .vdd(vdd), .A(_2618_), .B(_2937_), .C(_2948_), .Y(_2954_) );
AOI21X1 AOI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_2954_), .B(_2953_), .C(_2952_), .Y(_2955_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_2951_), .B(_2955_), .Y(_2956_) );
XNOR2X1 XNOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_2956_), .B(_2616_), .Y(H_22_) );
NAND3X1 NAND3X1_572 ( .gnd(gnd), .vdd(vdd), .A(_2952_), .B(_2954_), .C(_2953_), .Y(_2957_) );
OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_2616_), .B(_2955_), .C(_2957_), .Y(_2958_) );
OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_2911_), .B(_2621_), .C(_2914_), .Y(_2960_) );
OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2624_), .B(_2893_), .C(_2897_), .Y(_2961_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_2876_), .B(_2878_), .Y(_2962_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_2846_), .B(_2860_), .Y(_2963_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_2824_), .B(_2837_), .Y(_2964_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_2803_), .B(_2816_), .Y(_2965_) );
OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_2634_), .B(_2788_), .C(_2791_), .Y(_2966_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(_2786_), .Y(_2967_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .Y(_2968_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_2766_), .B(_2768_), .Y(_2969_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_2742_), .B(_2744_), .Y(_2971_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_2720_), .B(_2722_), .Y(_2972_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(_2972_), .Y(_2973_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_2698_), .B(_2700_), .Y(_2974_) );
OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_2676_), .B(_2643_), .C(_2678_), .Y(_2975_) );
OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .B(_2646_), .C(_2656_), .Y(_2976_) );
OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(W_12_), .B(W_13_), .C(W_14_), .Y(_2977_) );
XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(W_11_), .B(W_15_), .Y(_2978_) );
XNOR2X1 XNOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_2978_), .B(_2977_), .Y(_2979_) );
XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1551_), .B(W_31_), .Y(_2980_) );
XNOR2X1 XNOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_2980_), .B(_2979_), .Y(_2982_) );
XNOR2X1 XNOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_2653_), .B(_2982_), .Y(_2983_) );
XNOR2X1 XNOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_2983_), .B(_1360_), .Y(_2984_) );
XNOR2X1 XNOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1559_), .B(bloque_datos[15]), .Y(_2985_) );
XNOR2X1 XNOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_2984_), .B(_2985_), .Y(_2986_) );
XNOR2X1 XNOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_2986_), .B(_2976_), .Y(_2987_) );
XOR2X1 XOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_2987_), .B(_1566_), .Y(_2988_) );
NAND3X1 NAND3X1_573 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[14]), .B(_2664_), .C(_2668_), .Y(_2989_) );
XNOR2X1 XNOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .B(bloque_datos[31]), .Y(_2990_) );
XNOR2X1 XNOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_2990_), .B(_2989_), .Y(_2991_) );
XNOR2X1 XNOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_2988_), .B(_2991_), .Y(_2993_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_2975_), .B(_2993_), .Y(_2994_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(_2994_), .Y(_2995_) );
OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2673_), .B(_2683_), .C(_2993_), .Y(_2996_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_2996_), .B(_2995_), .Y(_2997_) );
AOI21X1 AOI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_3540_), .B(_3543_), .C(_2997_), .Y(_2998_) );
AOI21X1 AOI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_2996_), .B(_2995_), .C(_1587_), .Y(_2999_) );
XOR2X1 XOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1386_), .B(bloque_datos[47]), .Y(_3000_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(_3000_), .Y(_3001_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_3001_), .B(_2687_), .Y(_3002_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_2687_), .B(_3001_), .Y(_3004_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_3004_), .B(_3002_), .Y(_3005_) );
OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_2998_), .B(_2999_), .C(_3005_), .Y(_3006_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_2999_), .B(_2998_), .Y(_3007_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(_3007_), .Y(_3008_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_3005_), .B(_3008_), .Y(_3009_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(_3009_), .Y(_3010_) );
NAND3X1 NAND3X1_574 ( .gnd(gnd), .vdd(vdd), .A(_2974_), .B(_3006_), .C(_3010_), .Y(_3011_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(_2974_), .Y(_3012_) );
INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(_3006_), .Y(_3013_) );
OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_3009_), .B(_3013_), .C(_3012_), .Y(_3015_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_3557_), .B(_3553_), .Y(_3016_) );
XNOR2X1 XNOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .B(_3016_), .Y(_3017_) );
INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(_3017_), .Y(_3018_) );
AOI21X1 AOI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_3015_), .B(_3011_), .C(_3018_), .Y(_3019_) );
NAND3X1 NAND3X1_575 ( .gnd(gnd), .vdd(vdd), .A(_3012_), .B(_3006_), .C(_3010_), .Y(_3020_) );
OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_3009_), .B(_3013_), .C(_2974_), .Y(_3021_) );
AOI21X1 AOI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_3021_), .B(_3020_), .C(_3017_), .Y(_3022_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(_3022_), .Y(_3023_) );
XOR2X1 XOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_2708_), .B(bloque_datos[63]), .Y(_3024_) );
INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(_3024_), .Y(_3026_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_3026_), .B(_3023_), .Y(_3027_) );
OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(_3022_), .C(_3024_), .Y(_3028_) );
NAND3X1 NAND3X1_576 ( .gnd(gnd), .vdd(vdd), .A(_2973_), .B(_3028_), .C(_3027_), .Y(_3029_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_3023_), .B(_3026_), .Y(_3030_) );
INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(_3028_), .Y(_3031_) );
OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_3030_), .B(_3031_), .C(_2972_), .Y(_3032_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_3029_), .B(_3032_), .Y(_3033_) );
OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_3571_), .B(_3565_), .C(_3033_), .Y(_3034_) );
NAND3X1 NAND3X1_577 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .B(_3029_), .C(_3032_), .Y(_3035_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_3035_), .B(_3034_), .Y(_3037_) );
XOR2X1 XOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(bloque_datos[79]), .Y(_3038_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .B(_3038_), .Y(_3039_) );
INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .Y(_3040_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .B(_3038_), .Y(_3041_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_3041_), .B(_3040_), .Y(_3042_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_3042_), .B(_3037_), .Y(_3043_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_3037_), .B(_3042_), .Y(_3044_) );
NAND3X1 NAND3X1_578 ( .gnd(gnd), .vdd(vdd), .A(_2971_), .B(_3043_), .C(_3044_), .Y(_3045_) );
INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(_2971_), .Y(_3046_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_3037_), .B(_3042_), .Y(_3048_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_3042_), .B(_3037_), .Y(_3049_) );
OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_3048_), .B(_3049_), .C(_3046_), .Y(_3050_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(_1646_), .Y(_3051_) );
OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_3577_), .B(_3579_), .C(_1418_), .Y(_3052_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3051_), .B(_3052_), .C(_3050_), .D(_3045_), .Y(_3053_) );
NAND3X1 NAND3X1_579 ( .gnd(gnd), .vdd(vdd), .A(_3046_), .B(_3043_), .C(_3044_), .Y(_3054_) );
OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_3048_), .B(_3049_), .C(_2971_), .Y(_3055_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_3052_), .B(_3051_), .Y(_3056_) );
AOI21X1 AOI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .B(_3054_), .C(_3056_), .Y(_3057_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_3057_), .B(_3053_), .Y(_3059_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[95]), .B(_2754_), .Y(_3060_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[95]), .B(_2754_), .Y(_3061_) );
INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(_3061_), .Y(_3062_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_3060_), .B(_3062_), .Y(_3063_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_3063_), .B(_3059_), .Y(_3064_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_3059_), .B(_3063_), .Y(_3065_) );
NAND3X1 NAND3X1_580 ( .gnd(gnd), .vdd(vdd), .A(_2969_), .B(_3064_), .C(_3065_), .Y(_3066_) );
INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(_2969_), .Y(_3067_) );
INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(_3064_), .Y(_3068_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_3063_), .B(_3059_), .Y(_3070_) );
OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_3068_), .B(_3070_), .C(_3067_), .Y(_3071_) );
NAND3X1 NAND3X1_581 ( .gnd(gnd), .vdd(vdd), .A(_2968_), .B(_3066_), .C(_3071_), .Y(_3072_) );
NAND3X1 NAND3X1_582 ( .gnd(gnd), .vdd(vdd), .A(_3067_), .B(_3064_), .C(_3065_), .Y(_3073_) );
OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_3068_), .B(_3070_), .C(_2969_), .Y(_3074_) );
NAND3X1 NAND3X1_583 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .B(_3073_), .C(_3074_), .Y(_3075_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_3075_), .B(_3072_), .Y(_3076_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_2967_), .B(_3076_), .Y(_3077_) );
NAND3X1 NAND3X1_584 ( .gnd(gnd), .vdd(vdd), .A(_2786_), .B(_3075_), .C(_3072_), .Y(_3078_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_3078_), .B(_3077_), .Y(_3079_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_2966_), .B(_3079_), .Y(_3081_) );
INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(_2966_), .Y(_3082_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_3077_), .B(_3078_), .Y(_3083_) );
AOI21X1 AOI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_3082_), .B(_3083_), .C(_1536_), .Y(_3084_) );
XOR2X1 XOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_3603_), .B(W_143_), .Y(_3085_) );
NAND3X1 NAND3X1_585 ( .gnd(gnd), .vdd(vdd), .A(_3081_), .B(_3085_), .C(_3084_), .Y(_3086_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_3082_), .B(_3083_), .Y(_3087_) );
OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_3079_), .B(_2966_), .C(_1679_), .Y(_3088_) );
INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(_3085_), .Y(_3089_) );
OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_3087_), .B(_3088_), .C(_3089_), .Y(_3090_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_3090_), .B(_3086_), .Y(_3092_) );
XOR2X1 XOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_2798_), .Y(_3093_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_2965_), .B(_3093_), .Y(_3094_) );
INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(_2965_), .Y(_3095_) );
XNOR2X1 XNOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_2798_), .Y(_3096_) );
AOI21X1 AOI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .B(_3096_), .C(_1444_), .Y(_3097_) );
XOR2X1 XOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_3610_), .B(W_159_), .Y(_3098_) );
NAND3X1 NAND3X1_586 ( .gnd(gnd), .vdd(vdd), .A(_3094_), .B(_3098_), .C(_3097_), .Y(_3099_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .B(_3096_), .Y(_3100_) );
OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_3093_), .B(_2965_), .C(_1532_), .Y(_3101_) );
INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(_3098_), .Y(_3103_) );
OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .B(_3100_), .C(_3103_), .Y(_3104_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_3099_), .B(_3104_), .Y(_3105_) );
XOR2X1 XOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .B(_2820_), .Y(_3106_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_2964_), .B(_3106_), .Y(_3107_) );
INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(_2964_), .Y(_3108_) );
XNOR2X1 XNOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .B(_2820_), .Y(_3109_) );
AOI21X1 AOI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_3108_), .B(_3109_), .C(_1463_), .Y(_3110_) );
XOR2X1 XOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(W_175_), .Y(_3111_) );
NAND3X1 NAND3X1_587 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .B(_3111_), .C(_3110_), .Y(_3112_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_3108_), .B(_3109_), .Y(_3114_) );
OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_3106_), .B(_2964_), .C(_1457_), .Y(_3115_) );
INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3116_) );
OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_3115_), .B(_3114_), .C(_3116_), .Y(_3117_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_3112_), .B(_3117_), .Y(_3118_) );
XOR2X1 XOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_3118_), .B(_2841_), .Y(_3119_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_2963_), .B(_3119_), .Y(_3120_) );
INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(_2963_), .Y(_3121_) );
XNOR2X1 XNOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_3118_), .B(_2841_), .Y(_3122_) );
AOI21X1 AOI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_3121_), .B(_3122_), .C(_1472_), .Y(_3123_) );
XOR2X1 XOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_3622_), .B(W_191_), .Y(_3125_) );
NAND3X1 NAND3X1_588 ( .gnd(gnd), .vdd(vdd), .A(_3120_), .B(_3125_), .C(_3123_), .Y(_3126_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_3121_), .B(_3122_), .Y(_3127_) );
OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_3119_), .B(_2963_), .C(_1528_), .Y(_3128_) );
INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(_3125_), .Y(_3129_) );
OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_3128_), .B(_3127_), .C(_3129_), .Y(_3130_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_3126_), .B(_3130_), .Y(_3131_) );
XOR2X1 XOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_3131_), .B(_2870_), .Y(_3132_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_2962_), .B(_3132_), .Y(_3133_) );
INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(_2962_), .Y(_3134_) );
XNOR2X1 XNOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_3131_), .B(_2870_), .Y(_3136_) );
AOI21X1 AOI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_3134_), .B(_3136_), .C(_1484_), .Y(_3137_) );
XOR2X1 XOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_3629_), .B(W_207_), .Y(_3138_) );
NAND3X1 NAND3X1_589 ( .gnd(gnd), .vdd(vdd), .A(_3133_), .B(_3138_), .C(_3137_), .Y(_3139_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_3134_), .B(_3136_), .Y(_3140_) );
OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_3132_), .B(_2962_), .C(_1760_), .Y(_3141_) );
INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(_3138_), .Y(_3142_) );
OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_3141_), .B(_3140_), .C(_3142_), .Y(_3143_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_3139_), .B(_3143_), .Y(_3144_) );
XOR2X1 XOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_3144_), .B(_2891_), .Y(_3145_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_2961_), .B(_3145_), .Y(_3147_) );
INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(_2961_), .Y(_3148_) );
XNOR2X1 XNOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_3144_), .B(_2891_), .Y(_3149_) );
AOI21X1 AOI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_3148_), .B(_3149_), .C(_1496_), .Y(_3150_) );
XOR2X1 XOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_3634_), .B(W_223_), .Y(_3151_) );
NAND3X1 NAND3X1_590 ( .gnd(gnd), .vdd(vdd), .A(_3147_), .B(_3151_), .C(_3150_), .Y(_3152_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_3148_), .B(_3149_), .Y(_3153_) );
OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_3145_), .B(_2961_), .C(_1495_), .Y(_3154_) );
INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(_3151_), .Y(_3155_) );
OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_3154_), .B(_3153_), .C(_3155_), .Y(_3156_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_3152_), .B(_3156_), .Y(_3158_) );
XOR2X1 XOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_3158_), .B(_2909_), .Y(_3159_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_2960_), .B(_3159_), .Y(_3160_) );
INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(_2960_), .Y(_3161_) );
XNOR2X1 XNOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_3158_), .B(_2909_), .Y(_3162_) );
AOI21X1 AOI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_3161_), .B(_3162_), .C(_1510_), .Y(_3163_) );
XOR2X1 XOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(W_239_), .Y(_3164_) );
NAND3X1 NAND3X1_591 ( .gnd(gnd), .vdd(vdd), .A(_3160_), .B(_3164_), .C(_3163_), .Y(_3165_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_3161_), .B(_3162_), .Y(_3166_) );
OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_3159_), .B(_2960_), .C(_1509_), .Y(_3167_) );
XNOR2X1 XNOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(W_239_), .Y(_3169_) );
OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_3167_), .B(_3166_), .C(_3169_), .Y(_3170_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_3165_), .B(_3170_), .Y(_3171_) );
XOR2X1 XOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_3171_), .B(_2921_), .Y(_3172_) );
OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_2936_), .B(_2940_), .C(_3172_), .Y(_3173_) );
AOI21X1 AOI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_2931_), .B(_2620_), .C(_2940_), .Y(_3174_) );
XNOR2X1 XNOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_3171_), .B(_2921_), .Y(_3175_) );
AOI21X1 AOI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_3174_), .B(_3175_), .C(_1835_), .Y(_3176_) );
NAND3X1 NAND3X1_592 ( .gnd(gnd), .vdd(vdd), .A(W_255_), .B(_3173_), .C(_3176_), .Y(_3177_) );
INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(W_255_), .Y(_3178_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_3174_), .B(_3175_), .Y(_3180_) );
OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_2941_), .B(_2933_), .C(_2926_), .Y(_3181_) );
OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_3172_), .B(_3181_), .C(_1522_), .Y(_3182_) );
OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_3182_), .B(_3180_), .C(_3178_), .Y(_3183_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_3177_), .B(_3183_), .Y(_3184_) );
XNOR2X1 XNOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_3184_), .B(_2953_), .Y(_3185_) );
XNOR2X1 XNOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .B(_3185_), .Y(H_23_) );
INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(_1779_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(W_0_), .B(W_16_), .Y(_1790_) );
INVX2 INVX2_50 ( .gnd(gnd), .vdd(vdd), .A(W_0_), .Y(_1801_) );
INVX2 INVX2_51 ( .gnd(gnd), .vdd(vdd), .A(W_16_), .Y(_1812_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1801_), .B(_1812_), .Y(_1823_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1790_), .B(_1823_), .Y(_1834_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1779_), .B(_1834_), .Y(_1845_) );
OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_1823_), .B(_1790_), .C(bloque_datos[0]), .Y(_1856_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1856_), .B(_1845_), .Y(_1867_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .B(bloque_datos[16]), .Y(_1877_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[16]), .B(_1867_), .Y(_1886_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1886_), .B(_1877_), .Y(_1896_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_1896_), .B(bloque_datos[32]), .Y(_1906_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[32]), .B(_1896_), .Y(_1917_) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1917_), .B(_1906_), .Y(_1928_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .B(bloque_datos[48]), .Y(_1939_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[48]), .B(_1928_), .Y(_1950_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(_1939_), .Y(_1961_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_1961_), .B(bloque_datos[64]), .Y(_1972_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[64]), .B(_1961_), .Y(_1983_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1983_), .B(_1972_), .Y(_1994_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_1994_), .B(bloque_datos[80]), .Y(_2005_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .B(_1994_), .Y(_2016_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_2016_), .B(_2005_), .Y(_2027_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_2027_), .B(W_128_), .Y(_2038_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(W_128_), .B(_2027_), .Y(_2049_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_2049_), .B(_2038_), .Y(_2060_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(W_144_), .Y(_2071_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(W_144_), .B(_2060_), .Y(_2082_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_2082_), .B(_2071_), .Y(_2093_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_2093_), .B(W_160_), .Y(_2104_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(W_160_), .B(_2093_), .Y(_2115_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_2115_), .B(_2104_), .Y(_2126_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_2126_), .B(W_176_), .Y(_2137_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(W_176_), .B(_2126_), .Y(_2148_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_2148_), .B(_2137_), .Y(_2159_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_2159_), .B(W_192_), .Y(_2170_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(W_192_), .B(_2159_), .Y(_2181_) );
NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_2181_), .B(_2170_), .Y(_2192_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_2192_), .B(W_208_), .Y(_2203_) );
NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(W_208_), .B(_2192_), .Y(_2214_) );
NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_2214_), .B(_2203_), .Y(_2225_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_2225_), .B(W_224_), .Y(_2236_) );
NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(W_224_), .B(_2225_), .Y(_2247_) );
NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_2247_), .B(_2236_), .Y(_2257_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(_2257_), .Y(_2268_) );
INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(W_241_), .Y(_2279_) );
INVX2 INVX2_52 ( .gnd(gnd), .vdd(vdd), .A(_2225_), .Y(_2290_) );
INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(W_225_), .Y(_2301_) );
INVX2 INVX2_53 ( .gnd(gnd), .vdd(vdd), .A(_2192_), .Y(_2312_) );
INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(W_209_), .Y(_2323_) );
INVX2 INVX2_54 ( .gnd(gnd), .vdd(vdd), .A(_2159_), .Y(_2334_) );
INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(W_193_), .Y(_2345_) );
INVX2 INVX2_55 ( .gnd(gnd), .vdd(vdd), .A(_2126_), .Y(_2356_) );
INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(W_177_), .Y(_2367_) );
INVX2 INVX2_56 ( .gnd(gnd), .vdd(vdd), .A(_2093_), .Y(_2378_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(W_160_), .B(_2378_), .Y(_2389_) );
INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(W_161_), .Y(_2400_) );
INVX2 INVX2_57 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .Y(_2411_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(W_144_), .B(_2411_), .Y(_2422_) );
INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(W_145_), .Y(_2433_) );
INVX2 INVX2_58 ( .gnd(gnd), .vdd(vdd), .A(_2027_), .Y(_2444_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(W_128_), .B(_2444_), .Y(_2455_) );
INVX1 INVX1_264 ( .gnd(gnd), .vdd(vdd), .A(W_129_), .Y(_2466_) );
INVX2 INVX2_59 ( .gnd(gnd), .vdd(vdd), .A(_1994_), .Y(_2477_) );
INVX1 INVX1_265 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[81]), .Y(_2488_) );
INVX1 INVX1_266 ( .gnd(gnd), .vdd(vdd), .A(_1961_), .Y(_2499_) );
INVX1 INVX1_267 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[65]), .Y(_2510_) );
INVX1 INVX1_268 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .Y(_2521_) );
INVX1 INVX1_269 ( .gnd(gnd), .vdd(vdd), .A(_1896_), .Y(_2532_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[32]), .B(_2532_), .Y(_2543_) );
INVX1 INVX1_270 ( .gnd(gnd), .vdd(vdd), .A(_2543_), .Y(_2554_) );
INVX1 INVX1_271 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .Y(_2565_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[16]), .B(_2565_), .Y(_2576_) );
INVX1 INVX1_272 ( .gnd(gnd), .vdd(vdd), .A(_2576_), .Y(_2587_) );
OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1823_), .B(_1790_), .C(_1779_), .Y(_2598_) );
INVX1 INVX1_273 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(_2609_) );
INVX2 INVX2_60 ( .gnd(gnd), .vdd(vdd), .A(W_17_), .Y(_2619_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(W_0_), .B(W_1_), .Y(_2630_) );
INVX1 INVX1_274 ( .gnd(gnd), .vdd(vdd), .A(_2630_), .Y(_2641_) );
NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(W_0_), .B(W_1_), .Y(_2652_) );
NAND3X1 NAND3X1_593 ( .gnd(gnd), .vdd(vdd), .A(_2619_), .B(_2652_), .C(_2641_), .Y(_2663_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(_2652_), .Y(_2674_) );
OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_2674_), .B(_2630_), .C(W_17_), .Y(_2685_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(W_0_), .B(_1812_), .C(_2663_), .D(_2685_), .Y(_2696_) );
NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(W_0_), .B(_1812_), .Y(_2707_) );
NAND3X1 NAND3X1_594 ( .gnd(gnd), .vdd(vdd), .A(W_17_), .B(_2652_), .C(_2641_), .Y(_2718_) );
OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_2674_), .B(_2630_), .C(_2619_), .Y(_2729_) );
AOI21X1 AOI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_2729_), .B(_2718_), .C(_2707_), .Y(_2740_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .B(_2740_), .Y(_2751_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_2609_), .B(_2751_), .Y(_2762_) );
INVX2 INVX2_61 ( .gnd(gnd), .vdd(vdd), .A(_2762_), .Y(_2773_) );
OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .B(_2740_), .C(_2609_), .Y(_2784_) );
NAND3X1 NAND3X1_595 ( .gnd(gnd), .vdd(vdd), .A(_2598_), .B(_2784_), .C(_2773_), .Y(_2795_) );
INVX1 INVX1_275 ( .gnd(gnd), .vdd(vdd), .A(_2598_), .Y(_2806_) );
INVX1 INVX1_276 ( .gnd(gnd), .vdd(vdd), .A(_2784_), .Y(_2817_) );
OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_2762_), .B(_2817_), .C(_2806_), .Y(_2828_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_2795_), .B(_2828_), .Y(_2839_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_2839_), .B(bloque_datos[17]), .Y(_2850_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .B(_2839_), .Y(_2861_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_2861_), .B(_2850_), .Y(_2872_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_2872_), .B(_2587_), .Y(_2883_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_2587_), .B(_2872_), .Y(_2894_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_2894_), .B(_2883_), .Y(_2905_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_2905_), .B(bloque_datos[33]), .Y(_2916_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[33]), .B(_2905_), .Y(_2927_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_2927_), .B(_2916_), .Y(_2938_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_2938_), .B(_2554_), .Y(_2949_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_2554_), .B(_2938_), .Y(_2959_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .B(_2949_), .Y(_2970_) );
NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[49]), .B(_2970_), .Y(_2981_) );
INVX2 INVX2_62 ( .gnd(gnd), .vdd(vdd), .A(_2981_), .Y(_2992_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[49]), .B(_2970_), .Y(_3003_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_3003_), .B(_2992_), .Y(_3014_) );
OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[48]), .B(_2521_), .C(_3014_), .Y(_3025_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[48]), .B(_2521_), .Y(_3036_) );
OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2992_), .B(_3003_), .C(_3036_), .Y(_3047_) );
NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_3047_), .B(_3025_), .Y(_3058_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_2510_), .B(_3058_), .Y(_3069_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_3025_), .B(_3047_), .Y(_3080_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[65]), .B(_3080_), .Y(_3091_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_3069_), .B(_3091_), .Y(_3102_) );
OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[64]), .B(_2499_), .C(_3102_), .Y(_3113_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[64]), .B(_2499_), .Y(_3124_) );
OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_3091_), .B(_3069_), .C(_3124_), .Y(_3135_) );
NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_3135_), .B(_3113_), .Y(_3146_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_2488_), .B(_3146_), .Y(_3157_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .B(_3135_), .Y(_3168_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[81]), .B(_3168_), .Y(_3179_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_3157_), .B(_3179_), .Y(_3186_) );
OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .B(_2477_), .C(_3186_), .Y(_3187_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .B(_2477_), .Y(_3188_) );
OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_3179_), .B(_3157_), .C(_3188_), .Y(_3189_) );
NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_3189_), .B(_3187_), .Y(_3190_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_2466_), .B(_3190_), .Y(_3191_) );
INVX1 INVX1_277 ( .gnd(gnd), .vdd(vdd), .A(_3191_), .Y(_3192_) );
NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_2466_), .B(_3190_), .Y(_3193_) );
NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_3193_), .B(_3192_), .Y(_3194_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_2455_), .B(_3194_), .Y(_3195_) );
INVX1 INVX1_278 ( .gnd(gnd), .vdd(vdd), .A(_3195_), .Y(_3196_) );
NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2455_), .B(_3194_), .Y(_3197_) );
NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_3197_), .B(_3196_), .Y(_3198_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_2433_), .B(_3198_), .Y(_3199_) );
INVX1 INVX1_279 ( .gnd(gnd), .vdd(vdd), .A(_3199_), .Y(_3200_) );
NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_2433_), .B(_3198_), .Y(_3201_) );
NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_3201_), .B(_3200_), .Y(_3202_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_2422_), .B(_3202_), .Y(_3203_) );
INVX2 INVX2_63 ( .gnd(gnd), .vdd(vdd), .A(_3203_), .Y(_3204_) );
NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2422_), .B(_3202_), .Y(_3205_) );
NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_3205_), .B(_3204_), .Y(_3206_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_2400_), .B(_3206_), .Y(_3207_) );
INVX1 INVX1_280 ( .gnd(gnd), .vdd(vdd), .A(_3207_), .Y(_3208_) );
NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2400_), .B(_3206_), .Y(_3209_) );
NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_3209_), .B(_3208_), .Y(_3210_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .B(_3210_), .Y(_3211_) );
INVX2 INVX2_64 ( .gnd(gnd), .vdd(vdd), .A(_3211_), .Y(_3212_) );
NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .B(_3210_), .Y(_3213_) );
NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_3212_), .Y(_3214_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_2367_), .B(_3214_), .Y(_3215_) );
INVX2 INVX2_65 ( .gnd(gnd), .vdd(vdd), .A(_3214_), .Y(_3216_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(W_177_), .B(_3216_), .Y(_3217_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .B(_3217_), .Y(_3218_) );
OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(W_176_), .B(_2356_), .C(_3218_), .Y(_3219_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(W_176_), .B(_2356_), .Y(_3220_) );
OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_3217_), .B(_3215_), .C(_3220_), .Y(_3221_) );
NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_3221_), .B(_3219_), .Y(_3222_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_2345_), .B(_3222_), .Y(_3223_) );
INVX2 INVX2_66 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .Y(_3224_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(W_193_), .B(_3224_), .Y(_3225_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_3223_), .B(_3225_), .Y(_3226_) );
OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(W_192_), .B(_2334_), .C(_3226_), .Y(_3227_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(W_192_), .B(_2334_), .Y(_3228_) );
OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_3225_), .B(_3223_), .C(_3228_), .Y(_3229_) );
NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_3229_), .B(_3227_), .Y(_3230_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_2323_), .B(_3230_), .Y(_3231_) );
INVX2 INVX2_67 ( .gnd(gnd), .vdd(vdd), .A(_3230_), .Y(_3232_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(W_209_), .B(_3232_), .Y(_3233_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_3231_), .B(_3233_), .Y(_3234_) );
OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(W_208_), .B(_2312_), .C(_3234_), .Y(_3235_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(W_208_), .B(_2312_), .Y(_3236_) );
OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_3233_), .B(_3231_), .C(_3236_), .Y(_3237_) );
NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_3237_), .B(_3235_), .Y(_3238_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_2301_), .B(_3238_), .Y(_3239_) );
INVX1 INVX1_281 ( .gnd(gnd), .vdd(vdd), .A(_3239_), .Y(_3240_) );
NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_2301_), .B(_3238_), .Y(_3241_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_3240_), .B(_3241_), .Y(_3242_) );
OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(W_224_), .B(_2290_), .C(_3242_), .Y(_3243_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(W_224_), .B(_2290_), .Y(_3244_) );
INVX1 INVX1_282 ( .gnd(gnd), .vdd(vdd), .A(_3242_), .Y(_3245_) );
NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_3244_), .B(_3245_), .Y(_3246_) );
NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_3243_), .B(_3246_), .Y(_3247_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_2279_), .B(_3247_), .Y(_3248_) );
INVX2 INVX2_68 ( .gnd(gnd), .vdd(vdd), .A(_3247_), .Y(_3249_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(W_241_), .B(_3249_), .Y(_3250_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_3248_), .B(_3250_), .Y(_3251_) );
OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(W_240_), .B(_2268_), .C(_3251_), .Y(_3252_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(W_240_), .B(_2268_), .Y(_3253_) );
OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_3250_), .B(_3248_), .C(_3253_), .Y(_3254_) );
NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_3254_), .B(_3252_), .Y(_3255_) );
INVX2 INVX2_69 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .Y(H_13_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_2268_), .B(W_240_), .Y(_3256_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_3253_), .B(_3256_), .Y(H_0_) );
INVX1 INVX1_283 ( .gnd(gnd), .vdd(vdd), .A(H_0_), .Y(H_12_) );
OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_3253_), .B(_3256_), .C(H_13_), .Y(_3257_) );
INVX1 INVX1_284 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .Y(_3258_) );
AOI21X1 AOI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_3251_), .B(H_0_), .C(_3258_), .Y(H_1_) );
INVX1 INVX1_285 ( .gnd(gnd), .vdd(vdd), .A(_3248_), .Y(_3259_) );
INVX1 INVX1_286 ( .gnd(gnd), .vdd(vdd), .A(W_242_), .Y(_3260_) );
INVX1 INVX1_287 ( .gnd(gnd), .vdd(vdd), .A(_3243_), .Y(_3261_) );
INVX1 INVX1_288 ( .gnd(gnd), .vdd(vdd), .A(W_226_), .Y(_3262_) );
INVX1 INVX1_289 ( .gnd(gnd), .vdd(vdd), .A(_3231_), .Y(_3263_) );
INVX1 INVX1_290 ( .gnd(gnd), .vdd(vdd), .A(W_210_), .Y(_3264_) );
INVX1 INVX1_291 ( .gnd(gnd), .vdd(vdd), .A(_3223_), .Y(_3265_) );
INVX1 INVX1_292 ( .gnd(gnd), .vdd(vdd), .A(W_194_), .Y(_3266_) );
INVX1 INVX1_293 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .Y(_3267_) );
INVX1 INVX1_294 ( .gnd(gnd), .vdd(vdd), .A(W_178_), .Y(_3268_) );
INVX1 INVX1_295 ( .gnd(gnd), .vdd(vdd), .A(W_162_), .Y(_3269_) );
INVX1 INVX1_296 ( .gnd(gnd), .vdd(vdd), .A(W_146_), .Y(_3270_) );
INVX1 INVX1_297 ( .gnd(gnd), .vdd(vdd), .A(W_130_), .Y(_3271_) );
NOR3X1 NOR3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_3188_), .B(_3157_), .C(_3179_), .Y(_3272_) );
NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[81]), .B(_3168_), .Y(_3273_) );
INVX1 INVX1_298 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[82]), .Y(_3274_) );
NOR3X1 NOR3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_3124_), .B(_3069_), .C(_3091_), .Y(_3275_) );
INVX1 INVX1_299 ( .gnd(gnd), .vdd(vdd), .A(_3069_), .Y(_3276_) );
INVX1 INVX1_300 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[66]), .Y(_3277_) );
INVX1 INVX1_301 ( .gnd(gnd), .vdd(vdd), .A(_3036_), .Y(_3278_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_3014_), .B(_3278_), .Y(_3279_) );
INVX1 INVX1_302 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[50]), .Y(_3280_) );
INVX1 INVX1_303 ( .gnd(gnd), .vdd(vdd), .A(_2916_), .Y(_3281_) );
INVX1 INVX1_304 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[34]), .Y(_3282_) );
INVX1 INVX1_305 ( .gnd(gnd), .vdd(vdd), .A(_2850_), .Y(_3283_) );
INVX1 INVX1_306 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .Y(_3284_) );
INVX2 INVX2_70 ( .gnd(gnd), .vdd(vdd), .A(_2795_), .Y(_3285_) );
INVX1 INVX1_307 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[2]), .Y(_3286_) );
INVX1 INVX1_308 ( .gnd(gnd), .vdd(vdd), .A(W_18_), .Y(_3287_) );
NAND3X1 NAND3X1_596 ( .gnd(gnd), .vdd(vdd), .A(W_0_), .B(W_1_), .C(W_2_), .Y(_3288_) );
INVX1 INVX1_309 ( .gnd(gnd), .vdd(vdd), .A(_3288_), .Y(_3289_) );
AOI21X1 AOI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(W_0_), .B(W_1_), .C(W_2_), .Y(_3290_) );
NOR3X1 NOR3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_3287_), .B(_3290_), .C(_3289_), .Y(_3291_) );
INVX2 INVX2_71 ( .gnd(gnd), .vdd(vdd), .A(_3290_), .Y(_3292_) );
AOI21X1 AOI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_3288_), .B(_3292_), .C(W_18_), .Y(_3293_) );
OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_3291_), .B(_3293_), .C(_2718_), .Y(_3294_) );
NOR3X1 NOR3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_2619_), .B(_2630_), .C(_2674_), .Y(_3295_) );
NAND3X1 NAND3X1_597 ( .gnd(gnd), .vdd(vdd), .A(W_18_), .B(_3288_), .C(_3292_), .Y(_3296_) );
OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_3289_), .B(_3290_), .C(_3287_), .Y(_3297_) );
NAND3X1 NAND3X1_598 ( .gnd(gnd), .vdd(vdd), .A(_3295_), .B(_3296_), .C(_3297_), .Y(_3298_) );
AOI21X1 AOI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_3298_), .B(_3294_), .C(_2696_), .Y(_3299_) );
NAND3X1 NAND3X1_599 ( .gnd(gnd), .vdd(vdd), .A(_2707_), .B(_2729_), .C(_2718_), .Y(_3300_) );
AOI21X1 AOI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_3296_), .B(_3297_), .C(_3295_), .Y(_3301_) );
NOR3X1 NOR3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_3293_), .B(_2718_), .C(_3291_), .Y(_3302_) );
NOR3X1 NOR3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_3300_), .B(_3301_), .C(_3302_), .Y(_3303_) );
NOR3X1 NOR3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_3286_), .B(_3299_), .C(_3303_), .Y(_3304_) );
OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_3303_), .B(_3299_), .C(_3286_), .Y(_3305_) );
INVX1 INVX1_310 ( .gnd(gnd), .vdd(vdd), .A(_3305_), .Y(_3306_) );
OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .B(_3304_), .C(_2773_), .Y(_3307_) );
INVX2 INVX2_72 ( .gnd(gnd), .vdd(vdd), .A(_3304_), .Y(_3308_) );
NAND3X1 NAND3X1_600 ( .gnd(gnd), .vdd(vdd), .A(_2762_), .B(_3305_), .C(_3308_), .Y(_3309_) );
AOI21X1 AOI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_3307_), .B(_3309_), .C(_3285_), .Y(_3310_) );
AOI21X1 AOI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_3305_), .B(_3308_), .C(_2762_), .Y(_3311_) );
NOR3X1 NOR3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_2773_), .B(_3304_), .C(_3306_), .Y(_3312_) );
NOR3X1 NOR3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_2795_), .C(_3311_), .Y(_3313_) );
NOR3X1 NOR3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_3284_), .B(_3310_), .C(_3313_), .Y(_3314_) );
OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_3311_), .B(_3312_), .C(_2795_), .Y(_3315_) );
NAND3X1 NAND3X1_601 ( .gnd(gnd), .vdd(vdd), .A(_3307_), .B(_3285_), .C(_3309_), .Y(_3316_) );
AOI21X1 AOI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_3316_), .B(_3315_), .C(bloque_datos[18]), .Y(_3317_) );
OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_3314_), .B(_3317_), .C(_3283_), .Y(_3318_) );
NAND3X1 NAND3X1_602 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .B(_3316_), .C(_3315_), .Y(_3319_) );
OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .B(_3310_), .C(_3284_), .Y(_3320_) );
NAND3X1 NAND3X1_603 ( .gnd(gnd), .vdd(vdd), .A(_2850_), .B(_3319_), .C(_3320_), .Y(_3321_) );
AOI21X1 AOI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_3321_), .B(_3318_), .C(_2883_), .Y(_3322_) );
OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[16]), .B(_2565_), .C(_2872_), .Y(_3323_) );
AOI21X1 AOI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_3319_), .B(_3320_), .C(_2850_), .Y(_3324_) );
NOR3X1 NOR3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_3283_), .B(_3317_), .C(_3314_), .Y(_3325_) );
NOR3X1 NOR3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_3323_), .B(_3324_), .C(_3325_), .Y(_3326_) );
NOR3X1 NOR3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_3282_), .B(_3322_), .C(_3326_), .Y(_3327_) );
OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_3326_), .B(_3322_), .C(_3282_), .Y(_3328_) );
INVX1 INVX1_311 ( .gnd(gnd), .vdd(vdd), .A(_3328_), .Y(_3329_) );
OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_3329_), .B(_3327_), .C(_3281_), .Y(_3330_) );
INVX2 INVX2_73 ( .gnd(gnd), .vdd(vdd), .A(_3327_), .Y(_3331_) );
NAND3X1 NAND3X1_604 ( .gnd(gnd), .vdd(vdd), .A(_2916_), .B(_3328_), .C(_3331_), .Y(_3332_) );
AOI21X1 AOI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_3332_), .C(_2949_), .Y(_3333_) );
OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[32]), .B(_2532_), .C(_2938_), .Y(_3334_) );
AOI21X1 AOI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_3328_), .B(_3331_), .C(_2916_), .Y(_3335_) );
NOR3X1 NOR3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_3281_), .B(_3327_), .C(_3329_), .Y(_3336_) );
NOR3X1 NOR3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(_3334_), .C(_3335_), .Y(_3337_) );
NOR3X1 NOR3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_3280_), .B(_3333_), .C(_3337_), .Y(_3338_) );
OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_3335_), .B(_3336_), .C(_3334_), .Y(_3339_) );
NAND3X1 NAND3X1_605 ( .gnd(gnd), .vdd(vdd), .A(_2949_), .B(_3330_), .C(_3332_), .Y(_3340_) );
AOI21X1 AOI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_3340_), .B(_3339_), .C(bloque_datos[50]), .Y(_3341_) );
OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_3338_), .B(_3341_), .C(_2981_), .Y(_3342_) );
NAND3X1 NAND3X1_606 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[50]), .B(_3340_), .C(_3339_), .Y(_3343_) );
OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_3337_), .B(_3333_), .C(_3280_), .Y(_3344_) );
NAND3X1 NAND3X1_607 ( .gnd(gnd), .vdd(vdd), .A(_2992_), .B(_3343_), .C(_3344_), .Y(_3345_) );
AOI21X1 AOI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_3345_), .B(_3342_), .C(_3279_), .Y(_3346_) );
AOI21X1 AOI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_3343_), .B(_3344_), .C(_2992_), .Y(_3347_) );
NOR3X1 NOR3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_2981_), .B(_3341_), .C(_3338_), .Y(_3348_) );
NOR3X1 NOR3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_3348_), .B(_3347_), .C(_3025_), .Y(_3349_) );
NOR3X1 NOR3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_3346_), .B(_3277_), .C(_3349_), .Y(_3350_) );
OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_3348_), .B(_3347_), .C(_3025_), .Y(_3351_) );
NAND3X1 NAND3X1_608 ( .gnd(gnd), .vdd(vdd), .A(_3342_), .B(_3345_), .C(_3279_), .Y(_3352_) );
AOI21X1 AOI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_3351_), .B(_3352_), .C(bloque_datos[66]), .Y(_3353_) );
OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_3350_), .B(_3353_), .C(_3276_), .Y(_3354_) );
NAND3X1 NAND3X1_609 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[66]), .B(_3351_), .C(_3352_), .Y(_3355_) );
OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_3349_), .B(_3346_), .C(_3277_), .Y(_3356_) );
NAND3X1 NAND3X1_610 ( .gnd(gnd), .vdd(vdd), .A(_3069_), .B(_3355_), .C(_3356_), .Y(_3357_) );
AOI21X1 AOI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_3357_), .B(_3354_), .C(_3275_), .Y(_3358_) );
AOI21X1 AOI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_3355_), .B(_3356_), .C(_3069_), .Y(_3359_) );
NOR3X1 NOR3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_3276_), .B(_3353_), .C(_3350_), .Y(_3360_) );
NOR3X1 NOR3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_3360_), .B(_3359_), .C(_3113_), .Y(_3361_) );
NOR3X1 NOR3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_3274_), .B(_3358_), .C(_3361_), .Y(_3362_) );
OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_3360_), .B(_3359_), .C(_3113_), .Y(_3363_) );
NAND3X1 NAND3X1_611 ( .gnd(gnd), .vdd(vdd), .A(_3275_), .B(_3357_), .C(_3354_), .Y(_3364_) );
AOI21X1 AOI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_3364_), .B(_3363_), .C(bloque_datos[82]), .Y(_3365_) );
OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_3362_), .B(_3365_), .C(_3273_), .Y(_3366_) );
NAND3X1 NAND3X1_612 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[82]), .B(_3364_), .C(_3363_), .Y(_3367_) );
OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_3361_), .B(_3358_), .C(_3274_), .Y(_3368_) );
NAND3X1 NAND3X1_613 ( .gnd(gnd), .vdd(vdd), .A(_3157_), .B(_3367_), .C(_3368_), .Y(_3369_) );
AOI21X1 AOI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_3366_), .C(_3272_), .Y(_3370_) );
AOI21X1 AOI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_3367_), .B(_3368_), .C(_3157_), .Y(_3371_) );
NOR3X1 NOR3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_3273_), .B(_3365_), .C(_3362_), .Y(_3372_) );
NOR3X1 NOR3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_3371_), .B(_3372_), .C(_3187_), .Y(_3373_) );
NOR3X1 NOR3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_3271_), .B(_3370_), .C(_3373_), .Y(_3374_) );
OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_3372_), .B(_3371_), .C(_3187_), .Y(_3375_) );
NAND3X1 NAND3X1_614 ( .gnd(gnd), .vdd(vdd), .A(_3272_), .B(_3369_), .C(_3366_), .Y(_3376_) );
AOI21X1 AOI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_3376_), .B(_3375_), .C(W_130_), .Y(_3377_) );
OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_3374_), .B(_3377_), .C(_3192_), .Y(_3378_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_3377_), .B(_3374_), .Y(_3379_) );
NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_3191_), .B(_3379_), .Y(_3380_) );
AOI21X1 AOI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_3378_), .B(_3380_), .C(_3195_), .Y(_3381_) );
NAND3X1 NAND3X1_615 ( .gnd(gnd), .vdd(vdd), .A(_3378_), .B(_3380_), .C(_3195_), .Y(_3382_) );
INVX1 INVX1_312 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .Y(_3383_) );
NOR3X1 NOR3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_3270_), .B(_3381_), .C(_3383_), .Y(_3384_) );
INVX1 INVX1_313 ( .gnd(gnd), .vdd(vdd), .A(_3381_), .Y(_3385_) );
AOI21X1 AOI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .B(_3385_), .C(W_146_), .Y(_3386_) );
OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_3384_), .B(_3386_), .C(_3200_), .Y(_3387_) );
INVX2 INVX2_74 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3388_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .B(_3384_), .Y(_3389_) );
NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_3199_), .B(_3389_), .Y(_3390_) );
INVX1 INVX1_314 ( .gnd(gnd), .vdd(vdd), .A(_3390_), .Y(_3391_) );
OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .B(_3388_), .C(_3204_), .Y(_3392_) );
INVX1 INVX1_315 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .Y(_3393_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_3391_), .Y(_3394_) );
NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_3203_), .B(_3394_), .Y(_3395_) );
INVX1 INVX1_316 ( .gnd(gnd), .vdd(vdd), .A(_3395_), .Y(_3396_) );
NOR3X1 NOR3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .B(_3269_), .C(_3396_), .Y(_3397_) );
AOI21X1 AOI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_3395_), .C(W_162_), .Y(_3398_) );
OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_3397_), .B(_3398_), .C(_3208_), .Y(_3399_) );
INVX1 INVX1_317 ( .gnd(gnd), .vdd(vdd), .A(_3399_), .Y(_3400_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_3398_), .B(_3397_), .Y(_3401_) );
NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_3207_), .B(_3401_), .Y(_3402_) );
INVX1 INVX1_318 ( .gnd(gnd), .vdd(vdd), .A(_3402_), .Y(_3403_) );
OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_3403_), .B(_3400_), .C(_3212_), .Y(_3404_) );
INVX1 INVX1_319 ( .gnd(gnd), .vdd(vdd), .A(_3404_), .Y(_3405_) );
NAND3X1 NAND3X1_616 ( .gnd(gnd), .vdd(vdd), .A(_3211_), .B(_3399_), .C(_3402_), .Y(_3406_) );
INVX1 INVX1_320 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .Y(_3407_) );
NOR3X1 NOR3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_3268_), .B(_3407_), .C(_3405_), .Y(_3408_) );
AOI21X1 AOI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .B(_3404_), .C(W_178_), .Y(_3409_) );
OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .B(_3409_), .C(_3267_), .Y(_3410_) );
INVX1 INVX1_321 ( .gnd(gnd), .vdd(vdd), .A(_3410_), .Y(_3411_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_3409_), .B(_3408_), .Y(_3412_) );
NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .B(_3412_), .Y(_3413_) );
INVX1 INVX1_322 ( .gnd(gnd), .vdd(vdd), .A(_3413_), .Y(_3414_) );
OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_3414_), .B(_3411_), .C(_3219_), .Y(_3415_) );
INVX1 INVX1_323 ( .gnd(gnd), .vdd(vdd), .A(_3415_), .Y(_3416_) );
INVX1 INVX1_324 ( .gnd(gnd), .vdd(vdd), .A(_3219_), .Y(_3417_) );
NAND3X1 NAND3X1_617 ( .gnd(gnd), .vdd(vdd), .A(_3417_), .B(_3410_), .C(_3413_), .Y(_3418_) );
INVX2 INVX2_75 ( .gnd(gnd), .vdd(vdd), .A(_3418_), .Y(_3419_) );
NOR3X1 NOR3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_3266_), .B(_3419_), .C(_3416_), .Y(_3420_) );
AOI21X1 AOI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_3418_), .B(_3415_), .C(W_194_), .Y(_3421_) );
OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_3420_), .B(_3421_), .C(_3265_), .Y(_3422_) );
INVX2 INVX2_76 ( .gnd(gnd), .vdd(vdd), .A(_3422_), .Y(_3423_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_3421_), .B(_3420_), .Y(_3424_) );
NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_3223_), .B(_3424_), .Y(_3425_) );
INVX1 INVX1_325 ( .gnd(gnd), .vdd(vdd), .A(_3425_), .Y(_3426_) );
OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_3426_), .B(_3423_), .C(_3227_), .Y(_3427_) );
INVX2 INVX2_77 ( .gnd(gnd), .vdd(vdd), .A(_3427_), .Y(_3428_) );
INVX1 INVX1_326 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .Y(_3429_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_3423_), .B(_3426_), .Y(_3430_) );
NAND2X1 NAND2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_3429_), .B(_3430_), .Y(_3431_) );
INVX2 INVX2_78 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .Y(_3432_) );
NOR3X1 NOR3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_3264_), .B(_3428_), .C(_3432_), .Y(_3433_) );
AOI21X1 AOI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_3427_), .B(_3431_), .C(W_210_), .Y(_3434_) );
OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .B(_3434_), .C(_3263_), .Y(_3435_) );
INVX1 INVX1_327 ( .gnd(gnd), .vdd(vdd), .A(_3435_), .Y(_3436_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_3428_), .B(_3432_), .Y(_3437_) );
NAND2X1 NAND2X1_325 ( .gnd(gnd), .vdd(vdd), .A(W_210_), .B(_3437_), .Y(_3438_) );
INVX1 INVX1_328 ( .gnd(gnd), .vdd(vdd), .A(_3434_), .Y(_3439_) );
NAND3X1 NAND3X1_618 ( .gnd(gnd), .vdd(vdd), .A(_3231_), .B(_3439_), .C(_3438_), .Y(_3440_) );
INVX1 INVX1_329 ( .gnd(gnd), .vdd(vdd), .A(_3440_), .Y(_3441_) );
OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_3441_), .B(_3436_), .C(_3235_), .Y(_3442_) );
INVX2 INVX2_79 ( .gnd(gnd), .vdd(vdd), .A(_3442_), .Y(_3443_) );
INVX1 INVX1_330 ( .gnd(gnd), .vdd(vdd), .A(_3235_), .Y(_3444_) );
NAND3X1 NAND3X1_619 ( .gnd(gnd), .vdd(vdd), .A(_3444_), .B(_3435_), .C(_3440_), .Y(_3445_) );
INVX2 INVX2_80 ( .gnd(gnd), .vdd(vdd), .A(_3445_), .Y(_3446_) );
NOR3X1 NOR3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_3262_), .B(_3446_), .C(_3443_), .Y(_3447_) );
OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_3443_), .B(_3446_), .C(_3262_), .Y(_3448_) );
INVX1 INVX1_331 ( .gnd(gnd), .vdd(vdd), .A(_3448_), .Y(_3449_) );
OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_3449_), .B(_3447_), .C(_3240_), .Y(_3450_) );
INVX2 INVX2_81 ( .gnd(gnd), .vdd(vdd), .A(_3447_), .Y(_3451_) );
NAND3X1 NAND3X1_620 ( .gnd(gnd), .vdd(vdd), .A(_3239_), .B(_3448_), .C(_3451_), .Y(_3452_) );
AOI21X1 AOI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_3450_), .B(_3452_), .C(_3261_), .Y(_3453_) );
NAND3X1 NAND3X1_621 ( .gnd(gnd), .vdd(vdd), .A(_3261_), .B(_3450_), .C(_3452_), .Y(_3454_) );
INVX1 INVX1_332 ( .gnd(gnd), .vdd(vdd), .A(_3454_), .Y(_3455_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_3453_), .B(_3455_), .Y(_3456_) );
INVX2 INVX2_82 ( .gnd(gnd), .vdd(vdd), .A(_3456_), .Y(_3457_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_3260_), .B(_3457_), .Y(_3458_) );
OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_3455_), .B(_3453_), .C(_3260_), .Y(_3459_) );
INVX1 INVX1_333 ( .gnd(gnd), .vdd(vdd), .A(_3459_), .Y(_3460_) );
OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_3458_), .B(_3460_), .C(_3259_), .Y(_3461_) );
INVX1 INVX1_334 ( .gnd(gnd), .vdd(vdd), .A(_3461_), .Y(_3462_) );
INVX1 INVX1_335 ( .gnd(gnd), .vdd(vdd), .A(_3458_), .Y(_3463_) );
NAND3X1 NAND3X1_622 ( .gnd(gnd), .vdd(vdd), .A(_3248_), .B(_3459_), .C(_3463_), .Y(_3464_) );
INVX1 INVX1_336 ( .gnd(gnd), .vdd(vdd), .A(_3464_), .Y(_3465_) );
OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_3465_), .B(_3462_), .C(_3252_), .Y(_3466_) );
INVX1 INVX1_337 ( .gnd(gnd), .vdd(vdd), .A(_3252_), .Y(_3467_) );
NAND3X1 NAND3X1_623 ( .gnd(gnd), .vdd(vdd), .A(_3467_), .B(_3461_), .C(_3464_), .Y(_3468_) );
NAND2X1 NAND2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_3468_), .B(_3466_), .Y(_3469_) );
INVX2 INVX2_83 ( .gnd(gnd), .vdd(vdd), .A(_3469_), .Y(H_14_) );
NAND2X1 NAND2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_3258_), .B(H_14_), .Y(_3470_) );
OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(H_0_), .C(_3469_), .Y(_3471_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_3470_), .B(_3471_), .Y(H_2_) );
OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_3462_), .B(_3252_), .C(_3464_), .Y(_3472_) );
INVX2 INVX2_84 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .Y(_3473_) );
NAND2X1 NAND2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_3452_), .B(_3454_), .Y(_3474_) );
INVX1 INVX1_338 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .Y(_3475_) );
OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_3436_), .B(_3235_), .C(_3440_), .Y(_3476_) );
OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_3423_), .B(_3227_), .C(_3425_), .Y(_3477_) );
INVX1 INVX1_339 ( .gnd(gnd), .vdd(vdd), .A(_3477_), .Y(_3478_) );
INVX2 INVX2_85 ( .gnd(gnd), .vdd(vdd), .A(_3420_), .Y(_3479_) );
OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_3411_), .B(_3219_), .C(_3413_), .Y(_3480_) );
OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_3400_), .B(_3212_), .C(_3402_), .Y(_3481_) );
INVX1 INVX1_340 ( .gnd(gnd), .vdd(vdd), .A(_3481_), .Y(_3482_) );
INVX2 INVX2_86 ( .gnd(gnd), .vdd(vdd), .A(_3397_), .Y(_3483_) );
OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_3204_), .B(_3388_), .C(_3390_), .Y(_3484_) );
INVX1 INVX1_341 ( .gnd(gnd), .vdd(vdd), .A(W_147_), .Y(_3485_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .B(_3380_), .Y(_3486_) );
INVX1 INVX1_342 ( .gnd(gnd), .vdd(vdd), .A(W_131_), .Y(_3487_) );
OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_3187_), .B(_3371_), .C(_3369_), .Y(_3488_) );
INVX1 INVX1_343 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[83]), .Y(_3489_) );
OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .B(_3359_), .C(_3357_), .Y(_3490_) );
INVX2 INVX2_87 ( .gnd(gnd), .vdd(vdd), .A(_3490_), .Y(_3491_) );
INVX1 INVX1_344 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[67]), .Y(_3492_) );
OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_3025_), .B(_3347_), .C(_3345_), .Y(_3493_) );
INVX1 INVX1_345 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[51]), .Y(_3494_) );
OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_3335_), .B(_3334_), .C(_3332_), .Y(_3495_) );
INVX1 INVX1_346 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[35]), .Y(_3496_) );
INVX1 INVX1_347 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[19]), .Y(_3497_) );
AOI21X1 AOI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_3307_), .B(_3285_), .C(_3312_), .Y(_3498_) );
INVX1 INVX1_348 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[3]), .Y(_3499_) );
AOI21X1 AOI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .B(_3294_), .C(_3302_), .Y(_3500_) );
INVX1 INVX1_349 ( .gnd(gnd), .vdd(vdd), .A(W_19_), .Y(_3501_) );
INVX2 INVX2_88 ( .gnd(gnd), .vdd(vdd), .A(W_3_), .Y(_3502_) );
NAND2X1 NAND2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_3502_), .B(_3288_), .Y(_3503_) );
INVX1 INVX1_350 ( .gnd(gnd), .vdd(vdd), .A(_3503_), .Y(_3504_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_3502_), .B(_3288_), .Y(_3505_) );
NOR3X1 NOR3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_3501_), .B(_3505_), .C(_3504_), .Y(_3506_) );
INVX2 INVX2_89 ( .gnd(gnd), .vdd(vdd), .A(_3505_), .Y(_3507_) );
AOI21X1 AOI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_3503_), .B(_3507_), .C(W_19_), .Y(_3508_) );
OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_3506_), .C(_3291_), .Y(_3509_) );
NAND3X1 NAND3X1_624 ( .gnd(gnd), .vdd(vdd), .A(W_19_), .B(_3503_), .C(_3507_), .Y(_3510_) );
OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_3504_), .B(_3505_), .C(_3501_), .Y(_3511_) );
NAND3X1 NAND3X1_625 ( .gnd(gnd), .vdd(vdd), .A(_3296_), .B(_3511_), .C(_3510_), .Y(_3512_) );
NAND2X1 NAND2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_3512_), .B(_3509_), .Y(_3513_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_3500_), .B(_3513_), .Y(_3514_) );
OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_3301_), .B(_3300_), .C(_3298_), .Y(_3515_) );
AOI21X1 AOI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_3512_), .B(_3509_), .C(_3515_), .Y(_3516_) );
NOR3X1 NOR3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_3499_), .B(_3516_), .C(_3514_), .Y(_3517_) );
INVX1 INVX1_351 ( .gnd(gnd), .vdd(vdd), .A(_3517_), .Y(_3518_) );
OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_3514_), .B(_3516_), .C(_3499_), .Y(_3519_) );
AOI21X1 AOI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_3519_), .B(_3518_), .C(_3308_), .Y(_3520_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_3513_), .B(_3500_), .Y(_3521_) );
INVX1 INVX1_352 ( .gnd(gnd), .vdd(vdd), .A(_3516_), .Y(_3522_) );
AOI21X1 AOI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_3522_), .B(_3521_), .C(bloque_datos[3]), .Y(_3523_) );
NOR3X1 NOR3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_3517_), .B(_3304_), .C(_3523_), .Y(_3524_) );
NOR3X1 NOR3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_3524_), .C(_3520_), .Y(_3525_) );
OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_3311_), .B(_2795_), .C(_3309_), .Y(_3526_) );
OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_3523_), .B(_3517_), .C(_3304_), .Y(_3527_) );
NAND3X1 NAND3X1_626 ( .gnd(gnd), .vdd(vdd), .A(_3308_), .B(_3519_), .C(_3518_), .Y(_3528_) );
AOI21X1 AOI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_3527_), .B(_3528_), .C(_3526_), .Y(_3529_) );
OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_3525_), .B(_3529_), .C(_3497_), .Y(_3530_) );
NAND3X1 NAND3X1_627 ( .gnd(gnd), .vdd(vdd), .A(_3526_), .B(_3527_), .C(_3528_), .Y(_3531_) );
OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_3520_), .B(_3524_), .C(_3498_), .Y(_3532_) );
NAND3X1 NAND3X1_628 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[19]), .B(_3531_), .C(_3532_), .Y(_3533_) );
NAND3X1 NAND3X1_629 ( .gnd(gnd), .vdd(vdd), .A(_3319_), .B(_3533_), .C(_3530_), .Y(_3534_) );
NAND3X1 NAND3X1_630 ( .gnd(gnd), .vdd(vdd), .A(_3497_), .B(_3531_), .C(_3532_), .Y(_3535_) );
OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_3525_), .B(_3529_), .C(bloque_datos[19]), .Y(_3536_) );
NAND3X1 NAND3X1_631 ( .gnd(gnd), .vdd(vdd), .A(_3314_), .B(_3535_), .C(_3536_), .Y(_3537_) );
NAND2X1 NAND2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_3534_), .B(_3537_), .Y(_3538_) );
INVX1 INVX1_353 ( .gnd(gnd), .vdd(vdd), .A(_3538_), .Y(_3539_) );
OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_3325_), .B(_3326_), .C(_3539_), .Y(_3540_) );
OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_3324_), .B(_3323_), .C(_3321_), .Y(_3541_) );
INVX2 INVX2_90 ( .gnd(gnd), .vdd(vdd), .A(_3541_), .Y(_3542_) );
NAND2X1 NAND2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_3542_), .B(_3538_), .Y(_3543_) );
NAND3X1 NAND3X1_632 ( .gnd(gnd), .vdd(vdd), .A(_3496_), .B(_3543_), .C(_3540_), .Y(_3544_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_3542_), .B(_3538_), .Y(_3545_) );
INVX1 INVX1_354 ( .gnd(gnd), .vdd(vdd), .A(_3543_), .Y(_3546_) );
OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_3546_), .B(_3545_), .C(bloque_datos[35]), .Y(_3547_) );
AOI21X1 AOI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_3544_), .B(_3547_), .C(_3327_), .Y(_3548_) );
INVX1 INVX1_355 ( .gnd(gnd), .vdd(vdd), .A(_3548_), .Y(_3549_) );
NAND2X1 NAND2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_3544_), .B(_3547_), .Y(_3550_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_3550_), .B(_3331_), .Y(_3551_) );
NAND3X1 NAND3X1_633 ( .gnd(gnd), .vdd(vdd), .A(_3495_), .B(_3549_), .C(_3551_), .Y(_3552_) );
INVX2 INVX2_91 ( .gnd(gnd), .vdd(vdd), .A(_3552_), .Y(_3553_) );
INVX1 INVX1_356 ( .gnd(gnd), .vdd(vdd), .A(_3495_), .Y(_3554_) );
NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_3331_), .B(_3550_), .Y(_3555_) );
OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_3555_), .B(_3548_), .C(_3554_), .Y(_3556_) );
INVX2 INVX2_92 ( .gnd(gnd), .vdd(vdd), .A(_3556_), .Y(_3557_) );
OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .B(_3557_), .C(_3494_), .Y(_3558_) );
NAND3X1 NAND3X1_634 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[51]), .B(_3556_), .C(_3552_), .Y(_3559_) );
NAND3X1 NAND3X1_635 ( .gnd(gnd), .vdd(vdd), .A(_3343_), .B(_3559_), .C(_3558_), .Y(_3560_) );
NAND3X1 NAND3X1_636 ( .gnd(gnd), .vdd(vdd), .A(_3494_), .B(_3556_), .C(_3552_), .Y(_3561_) );
OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .B(_3557_), .C(bloque_datos[51]), .Y(_3562_) );
NAND3X1 NAND3X1_637 ( .gnd(gnd), .vdd(vdd), .A(_3338_), .B(_3561_), .C(_3562_), .Y(_3563_) );
NAND3X1 NAND3X1_638 ( .gnd(gnd), .vdd(vdd), .A(_3493_), .B(_3560_), .C(_3563_), .Y(_3564_) );
AOI21X1 AOI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_3560_), .B(_3563_), .C(_3493_), .Y(_3565_) );
INVX1 INVX1_357 ( .gnd(gnd), .vdd(vdd), .A(_3565_), .Y(_3566_) );
NAND3X1 NAND3X1_639 ( .gnd(gnd), .vdd(vdd), .A(_3492_), .B(_3564_), .C(_3566_), .Y(_3567_) );
INVX1 INVX1_358 ( .gnd(gnd), .vdd(vdd), .A(_3493_), .Y(_3568_) );
AOI21X1 AOI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_3561_), .B(_3562_), .C(_3338_), .Y(_3569_) );
AOI21X1 AOI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_3559_), .B(_3558_), .C(_3343_), .Y(_3570_) );
NOR3X1 NOR3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_3569_), .B(_3568_), .C(_3570_), .Y(_3571_) );
OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_3571_), .B(_3565_), .C(bloque_datos[67]), .Y(_3572_) );
AOI21X1 AOI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_3572_), .B(_3567_), .C(_3350_), .Y(_3573_) );
OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_3571_), .B(_3565_), .C(_3492_), .Y(_3574_) );
NAND3X1 NAND3X1_640 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[67]), .B(_3564_), .C(_3566_), .Y(_3575_) );
AOI21X1 AOI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .B(_3575_), .C(_3355_), .Y(_3576_) );
NOR3X1 NOR3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_3573_), .B(_3491_), .C(_3576_), .Y(_3577_) );
OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_3573_), .B(_3576_), .C(_3491_), .Y(_3578_) );
INVX2 INVX2_93 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .Y(_3579_) );
OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_3579_), .B(_3577_), .C(_3489_), .Y(_3580_) );
INVX2 INVX2_94 ( .gnd(gnd), .vdd(vdd), .A(_3577_), .Y(_3581_) );
NAND3X1 NAND3X1_641 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[83]), .B(_3578_), .C(_3581_), .Y(_3582_) );
NAND3X1 NAND3X1_642 ( .gnd(gnd), .vdd(vdd), .A(_3367_), .B(_3580_), .C(_3582_), .Y(_3583_) );
NAND3X1 NAND3X1_643 ( .gnd(gnd), .vdd(vdd), .A(_3489_), .B(_3578_), .C(_3581_), .Y(_3584_) );
OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_3579_), .B(_3577_), .C(bloque_datos[83]), .Y(_3585_) );
NAND3X1 NAND3X1_644 ( .gnd(gnd), .vdd(vdd), .A(_3362_), .B(_3585_), .C(_3584_), .Y(_3586_) );
NAND3X1 NAND3X1_645 ( .gnd(gnd), .vdd(vdd), .A(_3488_), .B(_3583_), .C(_3586_), .Y(_3587_) );
AOI21X1 AOI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_3583_), .B(_3586_), .C(_3488_), .Y(_3588_) );
INVX1 INVX1_359 ( .gnd(gnd), .vdd(vdd), .A(_3588_), .Y(_3589_) );
NAND3X1 NAND3X1_646 ( .gnd(gnd), .vdd(vdd), .A(_3487_), .B(_3587_), .C(_3589_), .Y(_3590_) );
INVX2 INVX2_95 ( .gnd(gnd), .vdd(vdd), .A(_3587_), .Y(_3591_) );
OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_3591_), .B(_3588_), .C(W_131_), .Y(_3592_) );
AOI21X1 AOI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_3590_), .B(_3592_), .C(_3374_), .Y(_3593_) );
INVX1 INVX1_360 ( .gnd(gnd), .vdd(vdd), .A(_3374_), .Y(_3594_) );
OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_3591_), .B(_3588_), .C(_3487_), .Y(_3595_) );
NAND3X1 NAND3X1_647 ( .gnd(gnd), .vdd(vdd), .A(W_131_), .B(_3587_), .C(_3589_), .Y(_3596_) );
AOI21X1 AOI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_3596_), .B(_3595_), .C(_3594_), .Y(_3597_) );
OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_3593_), .B(_3597_), .C(_3486_), .Y(_3598_) );
NAND2X1 NAND2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_3380_), .B(_3382_), .Y(_3599_) );
NAND3X1 NAND3X1_648 ( .gnd(gnd), .vdd(vdd), .A(_3594_), .B(_3596_), .C(_3595_), .Y(_3600_) );
NAND3X1 NAND3X1_649 ( .gnd(gnd), .vdd(vdd), .A(_3374_), .B(_3590_), .C(_3592_), .Y(_3601_) );
NAND3X1 NAND3X1_650 ( .gnd(gnd), .vdd(vdd), .A(_3600_), .B(_3601_), .C(_3599_), .Y(_3602_) );
NAND2X1 NAND2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_3602_), .B(_3598_), .Y(_3603_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_3603_), .B(_3485_), .Y(_3604_) );
NAND2X1 NAND2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_3485_), .B(_3603_), .Y(_3605_) );
NAND2X1 NAND2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_3605_), .B(_3604_), .Y(_3606_) );
XNOR2X1 XNOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_3606_), .B(_3384_), .Y(_3607_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_3607_), .B(_3484_), .Y(_3608_) );
NAND2X1 NAND2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_3484_), .B(_3607_), .Y(_3609_) );
NAND2X1 NAND2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_3609_), .B(_3608_), .Y(_3610_) );
XOR2X1 XOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_3610_), .B(W_163_), .Y(_3611_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_3611_), .B(_3483_), .Y(_3612_) );
NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_3483_), .B(_3611_), .Y(_3613_) );
OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_3612_), .B(_3613_), .C(_3482_), .Y(_3614_) );
NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_3613_), .B(_3612_), .Y(_3615_) );
NAND2X1 NAND2X1_340 ( .gnd(gnd), .vdd(vdd), .A(_3481_), .B(_3615_), .Y(_3616_) );
NAND2X1 NAND2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_3614_), .B(_3616_), .Y(_3617_) );
XOR2X1 XOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(W_179_), .Y(_3618_) );
XNOR2X1 XNOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_3618_), .B(_3408_), .Y(_3619_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_3619_), .B(_3480_), .Y(_3620_) );
OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_3419_), .B(_3414_), .C(_3619_), .Y(_3621_) );
NAND2X1 NAND2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_3621_), .B(_3620_), .Y(_3622_) );
XOR2X1 XOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_3622_), .B(W_195_), .Y(_3623_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_3623_), .B(_3479_), .Y(_3624_) );
NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_3479_), .B(_3623_), .Y(_3625_) );
OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_3624_), .B(_3625_), .C(_3478_), .Y(_3626_) );
NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_3625_), .B(_3624_), .Y(_3627_) );
NAND2X1 NAND2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_3477_), .B(_3627_), .Y(_3628_) );
NAND2X1 NAND2X1_344 ( .gnd(gnd), .vdd(vdd), .A(_3626_), .B(_3628_), .Y(_3629_) );
XOR2X1 XOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_3629_), .B(W_211_), .Y(_3630_) );
XNOR2X1 XNOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_3630_), .B(_3433_), .Y(_3631_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_3476_), .B(_3631_), .Y(_3632_) );
OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_3446_), .B(_3441_), .C(_3631_), .Y(_3633_) );
NAND2X1 NAND2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_3632_), .B(_3633_), .Y(_3634_) );
XOR2X1 XOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_3634_), .B(W_227_), .Y(_3635_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_3635_), .B(_3451_), .Y(_3636_) );
NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .B(_3635_), .Y(_3637_) );
OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_3636_), .B(_3637_), .C(_3475_), .Y(_3638_) );
NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_3637_), .B(_3636_), .Y(_3639_) );
NAND2X1 NAND2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .B(_3639_), .Y(_3640_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_3638_), .B(_3640_), .Y(_3641_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_3641_), .B(W_243_), .Y(_3642_) );
NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(W_243_), .B(_3641_), .Y(_3643_) );
OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_3642_), .B(_3643_), .C(_3463_), .Y(_3644_) );
NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_3643_), .B(_3642_), .Y(_3645_) );
NAND2X1 NAND2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_3458_), .B(_3645_), .Y(_3646_) );
NAND2X1 NAND2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3646_), .Y(_3647_) );
XNOR2X1 XNOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_3647_), .B(_3473_), .Y(H_15_) );
NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(H_15_), .B(_3470_), .Y(_3648_) );
INVX1 INVX1_361 ( .gnd(gnd), .vdd(vdd), .A(_3648_), .Y(_3649_) );
OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_3469_), .B(_3257_), .C(H_15_), .Y(_3650_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_3649_), .B(_3650_), .Y(H_3_) );
OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_3647_), .B(_3473_), .C(_3646_), .Y(_3651_) );
AOI21X1 AOI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .B(_3639_), .C(_3637_), .Y(_3652_) );
INVX2 INVX2_96 ( .gnd(gnd), .vdd(vdd), .A(_3652_), .Y(_3653_) );
INVX1 INVX1_362 ( .gnd(gnd), .vdd(vdd), .A(_3634_), .Y(_3654_) );
NAND2X1 NAND2X1_349 ( .gnd(gnd), .vdd(vdd), .A(W_227_), .B(_3654_), .Y(_3655_) );
INVX1 INVX1_363 ( .gnd(gnd), .vdd(vdd), .A(_3655_), .Y(_3656_) );
NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_3438_), .B(_3630_), .Y(_3657_) );
AOI21X1 AOI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_3631_), .B(_3476_), .C(_3657_), .Y(_3658_) );
INVX2 INVX2_97 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .Y(_3659_) );
INVX1 INVX1_364 ( .gnd(gnd), .vdd(vdd), .A(_3629_), .Y(_3660_) );
NAND2X1 NAND2X1_350 ( .gnd(gnd), .vdd(vdd), .A(W_211_), .B(_3660_), .Y(_3661_) );
INVX2 INVX2_98 ( .gnd(gnd), .vdd(vdd), .A(_3661_), .Y(_3662_) );
OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_3479_), .B(_3623_), .C(_3628_), .Y(_3663_) );
INVX1 INVX1_365 ( .gnd(gnd), .vdd(vdd), .A(_3622_), .Y(_3664_) );
NAND2X1 NAND2X1_351 ( .gnd(gnd), .vdd(vdd), .A(W_195_), .B(_3664_), .Y(_3665_) );
INVX2 INVX2_99 ( .gnd(gnd), .vdd(vdd), .A(_3665_), .Y(_3666_) );
INVX1 INVX1_366 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .Y(_3667_) );
OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_3667_), .B(_3618_), .C(_3621_), .Y(_3668_) );
INVX1 INVX1_367 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .Y(_3669_) );
NAND2X1 NAND2X1_352 ( .gnd(gnd), .vdd(vdd), .A(W_179_), .B(_3669_), .Y(_3670_) );
INVX1 INVX1_368 ( .gnd(gnd), .vdd(vdd), .A(_3670_), .Y(_3671_) );
OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_3483_), .B(_3611_), .C(_3616_), .Y(_3672_) );
INVX1 INVX1_369 ( .gnd(gnd), .vdd(vdd), .A(_3610_), .Y(_3673_) );
NAND2X1 NAND2X1_353 ( .gnd(gnd), .vdd(vdd), .A(W_163_), .B(_3673_), .Y(_3674_) );
INVX1 INVX1_370 ( .gnd(gnd), .vdd(vdd), .A(_3674_), .Y(_3675_) );
INVX1 INVX1_371 ( .gnd(gnd), .vdd(vdd), .A(_3384_), .Y(_3676_) );
OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_3676_), .B(_3606_), .C(_3609_), .Y(_3677_) );
INVX1 INVX1_372 ( .gnd(gnd), .vdd(vdd), .A(_3604_), .Y(_3678_) );
AOI21X1 AOI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_3600_), .B(_3599_), .C(_3597_), .Y(_3679_) );
INVX2 INVX2_100 ( .gnd(gnd), .vdd(vdd), .A(_3679_), .Y(_3680_) );
INVX1 INVX1_373 ( .gnd(gnd), .vdd(vdd), .A(W_132_), .Y(_3681_) );
NAND2X1 NAND2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_3586_), .B(_3587_), .Y(_3682_) );
INVX1 INVX1_374 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[84]), .Y(_3683_) );
INVX1 INVX1_375 ( .gnd(gnd), .vdd(vdd), .A(_3576_), .Y(_3684_) );
OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_3573_), .B(_3491_), .C(_3684_), .Y(_3685_) );
INVX1 INVX1_376 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[68]), .Y(_3686_) );
OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_3569_), .B(_3568_), .C(_3563_), .Y(_3687_) );
INVX1 INVX1_377 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[52]), .Y(_3688_) );
OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_3554_), .B(_3548_), .C(_3551_), .Y(_3689_) );
OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_3546_), .B(_3545_), .C(_3496_), .Y(_3690_) );
INVX1 INVX1_378 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[36]), .Y(_3691_) );
OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_3538_), .B(_3542_), .C(_3537_), .Y(_3692_) );
INVX1 INVX1_379 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[20]), .Y(_3693_) );
AOI21X1 AOI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_3526_), .B(_3528_), .C(_3520_), .Y(_3694_) );
AOI21X1 AOI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_3511_), .B(_3510_), .C(_3296_), .Y(_3695_) );
AOI21X1 AOI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_3512_), .B(_3515_), .C(_3695_), .Y(_3696_) );
INVX1 INVX1_380 ( .gnd(gnd), .vdd(vdd), .A(W_20_), .Y(_3697_) );
INVX1 INVX1_381 ( .gnd(gnd), .vdd(vdd), .A(W_4_), .Y(_3698_) );
NOR3X1 NOR3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_3502_), .B(_3698_), .C(_3288_), .Y(_3699_) );
OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_3288_), .B(_3502_), .C(_3698_), .Y(_3700_) );
INVX1 INVX1_382 ( .gnd(gnd), .vdd(vdd), .A(_3700_), .Y(_3701_) );
NOR3X1 NOR3X1_91 ( .gnd(gnd), .vdd(vdd), .A(W_0_), .B(_3699_), .C(_3701_), .Y(_3702_) );
NAND2X1 NAND2X1_355 ( .gnd(gnd), .vdd(vdd), .A(W_4_), .B(_3505_), .Y(_3703_) );
AOI21X1 AOI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_3700_), .B(_3703_), .C(_1801_), .Y(_3704_) );
OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_3702_), .B(_3704_), .C(_3697_), .Y(_3705_) );
NAND3X1 NAND3X1_651 ( .gnd(gnd), .vdd(vdd), .A(_1801_), .B(_3700_), .C(_3703_), .Y(_3706_) );
OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_3701_), .B(_3699_), .C(W_0_), .Y(_3707_) );
NAND3X1 NAND3X1_652 ( .gnd(gnd), .vdd(vdd), .A(W_20_), .B(_3706_), .C(_3707_), .Y(_3708_) );
NAND3X1 NAND3X1_653 ( .gnd(gnd), .vdd(vdd), .A(_3511_), .B(_3708_), .C(_3705_), .Y(_3709_) );
NAND3X1 NAND3X1_654 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3706_), .C(_3707_), .Y(_3710_) );
OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_3702_), .B(_3704_), .C(W_20_), .Y(_3711_) );
NAND3X1 NAND3X1_655 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_3710_), .C(_3711_), .Y(_3712_) );
NAND3X1 NAND3X1_656 ( .gnd(gnd), .vdd(vdd), .A(_3696_), .B(_3709_), .C(_3712_), .Y(_3713_) );
NOR3X1 NOR3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3506_), .B(_3291_), .C(_3508_), .Y(_3714_) );
OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_3500_), .B(_3714_), .C(_3509_), .Y(_3715_) );
NAND3X1 NAND3X1_657 ( .gnd(gnd), .vdd(vdd), .A(_3511_), .B(_3710_), .C(_3711_), .Y(_3716_) );
NAND3X1 NAND3X1_658 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_3708_), .C(_3705_), .Y(_3717_) );
NAND3X1 NAND3X1_659 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(_3717_), .C(_3715_), .Y(_3718_) );
XNOR2X1 XNOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1834_), .B(W_8_), .Y(_3719_) );
INVX1 INVX1_383 ( .gnd(gnd), .vdd(vdd), .A(_3719_), .Y(_3720_) );
NAND3X1 NAND3X1_660 ( .gnd(gnd), .vdd(vdd), .A(_3720_), .B(_3713_), .C(_3718_), .Y(_3721_) );
AOI21X1 AOI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(_3717_), .C(_3715_), .Y(_3722_) );
AOI21X1 AOI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_3709_), .B(_3712_), .C(_3696_), .Y(_3723_) );
OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .B(_3723_), .C(_3719_), .Y(_3724_) );
NAND3X1 NAND3X1_661 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[4]), .B(_3721_), .C(_3724_), .Y(_3725_) );
INVX1 INVX1_384 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[4]), .Y(_3726_) );
NAND3X1 NAND3X1_662 ( .gnd(gnd), .vdd(vdd), .A(_3719_), .B(_3713_), .C(_3718_), .Y(_3727_) );
OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .B(_3723_), .C(_3720_), .Y(_3728_) );
NAND3X1 NAND3X1_663 ( .gnd(gnd), .vdd(vdd), .A(_3726_), .B(_3727_), .C(_3728_), .Y(_3729_) );
NAND3X1 NAND3X1_664 ( .gnd(gnd), .vdd(vdd), .A(_3519_), .B(_3725_), .C(_3729_), .Y(_3730_) );
AOI21X1 AOI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_3727_), .B(_3728_), .C(_3726_), .Y(_3731_) );
AOI21X1 AOI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_3721_), .B(_3724_), .C(bloque_datos[4]), .Y(_3732_) );
OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_3731_), .B(_3732_), .C(_3523_), .Y(_3733_) );
AOI21X1 AOI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .B(_3733_), .C(_3694_), .Y(_3734_) );
OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_3524_), .C(_3527_), .Y(_3735_) );
OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_3731_), .B(_3732_), .C(_3519_), .Y(_3736_) );
NAND3X1 NAND3X1_665 ( .gnd(gnd), .vdd(vdd), .A(_3523_), .B(_3725_), .C(_3729_), .Y(_3737_) );
AOI21X1 AOI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_3737_), .B(_3736_), .C(_3735_), .Y(_3738_) );
NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(W_24_), .B(W_8_), .Y(_3739_) );
INVX1 INVX1_385 ( .gnd(gnd), .vdd(vdd), .A(_3739_), .Y(_3740_) );
NAND2X1 NAND2X1_356 ( .gnd(gnd), .vdd(vdd), .A(W_24_), .B(W_8_), .Y(_3741_) );
NAND2X1 NAND2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_3741_), .B(_3740_), .Y(_3742_) );
XNOR2X1 XNOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .B(_3742_), .Y(_3743_) );
OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_3734_), .B(_3738_), .C(_3743_), .Y(_3744_) );
NAND3X1 NAND3X1_666 ( .gnd(gnd), .vdd(vdd), .A(_3737_), .B(_3735_), .C(_3736_), .Y(_3745_) );
NAND3X1 NAND3X1_667 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .B(_3733_), .C(_3694_), .Y(_3746_) );
INVX1 INVX1_386 ( .gnd(gnd), .vdd(vdd), .A(_3743_), .Y(_3747_) );
NAND3X1 NAND3X1_668 ( .gnd(gnd), .vdd(vdd), .A(_3747_), .B(_3745_), .C(_3746_), .Y(_3748_) );
AOI21X1 AOI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .B(_3744_), .C(_3693_), .Y(_3749_) );
NAND3X1 NAND3X1_669 ( .gnd(gnd), .vdd(vdd), .A(_3743_), .B(_3745_), .C(_3746_), .Y(_3750_) );
OAI21X1 OAI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_3734_), .B(_3738_), .C(_3747_), .Y(_3751_) );
AOI21X1 AOI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_3750_), .B(_3751_), .C(bloque_datos[20]), .Y(_3752_) );
OAI21X1 OAI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_3749_), .B(_3752_), .C(_3530_), .Y(_3753_) );
INVX1 INVX1_387 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .Y(_3754_) );
NAND3X1 NAND3X1_670 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[20]), .B(_3750_), .C(_3751_), .Y(_3755_) );
NAND3X1 NAND3X1_671 ( .gnd(gnd), .vdd(vdd), .A(_3693_), .B(_3748_), .C(_3744_), .Y(_3756_) );
NAND3X1 NAND3X1_672 ( .gnd(gnd), .vdd(vdd), .A(_3754_), .B(_3755_), .C(_3756_), .Y(_3757_) );
NAND3X1 NAND3X1_673 ( .gnd(gnd), .vdd(vdd), .A(_3692_), .B(_3757_), .C(_3753_), .Y(_3758_) );
INVX1 INVX1_388 ( .gnd(gnd), .vdd(vdd), .A(_3537_), .Y(_3759_) );
AOI21X1 AOI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_3541_), .B(_3534_), .C(_3759_), .Y(_3760_) );
NAND3X1 NAND3X1_674 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(_3755_), .C(_3756_), .Y(_3761_) );
OAI21X1 OAI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_3749_), .B(_3752_), .C(_3754_), .Y(_3762_) );
NAND3X1 NAND3X1_675 ( .gnd(gnd), .vdd(vdd), .A(_3760_), .B(_3761_), .C(_3762_), .Y(_3763_) );
INVX1 INVX1_389 ( .gnd(gnd), .vdd(vdd), .A(_3742_), .Y(_3764_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_3764_), .B(bloque_datos[8]), .Y(_3765_) );
NAND2X1 NAND2X1_358 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .B(_3764_), .Y(_3766_) );
NAND2X1 NAND2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_3766_), .B(_3765_), .Y(_3767_) );
INVX2 INVX2_101 ( .gnd(gnd), .vdd(vdd), .A(_3767_), .Y(_3768_) );
XNOR2X1 XNOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1896_), .B(_3768_), .Y(_3769_) );
INVX1 INVX1_390 ( .gnd(gnd), .vdd(vdd), .A(_3769_), .Y(_3770_) );
NAND3X1 NAND3X1_676 ( .gnd(gnd), .vdd(vdd), .A(_3770_), .B(_3758_), .C(_3763_), .Y(_3771_) );
AOI21X1 AOI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_3761_), .B(_3762_), .C(_3760_), .Y(_2_) );
AOI21X1 AOI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_3757_), .B(_3753_), .C(_3692_), .Y(_3_) );
OAI21X1 OAI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(_3_), .C(_3769_), .Y(_4_) );
AOI21X1 AOI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_3771_), .B(_4_), .C(_3691_), .Y(_5_) );
NAND3X1 NAND3X1_677 ( .gnd(gnd), .vdd(vdd), .A(_3769_), .B(_3758_), .C(_3763_), .Y(_6_) );
OAI21X1 OAI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(_3_), .C(_3770_), .Y(_7_) );
AOI21X1 AOI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_7_), .C(bloque_datos[36]), .Y(_8_) );
OAI21X1 OAI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_8_), .C(_3690_), .Y(_9_) );
INVX1 INVX1_391 ( .gnd(gnd), .vdd(vdd), .A(_3690_), .Y(_10_) );
NAND3X1 NAND3X1_678 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[36]), .B(_6_), .C(_7_), .Y(_11_) );
NAND3X1 NAND3X1_679 ( .gnd(gnd), .vdd(vdd), .A(_3691_), .B(_3771_), .C(_4_), .Y(_12_) );
NAND3X1 NAND3X1_680 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_11_), .C(_12_), .Y(_13_) );
NAND3X1 NAND3X1_681 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_3689_), .C(_9_), .Y(_14_) );
AOI21X1 AOI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_3495_), .B(_3549_), .C(_3555_), .Y(_15_) );
NAND3X1 NAND3X1_682 ( .gnd(gnd), .vdd(vdd), .A(_3690_), .B(_11_), .C(_12_), .Y(_16_) );
OAI21X1 OAI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_8_), .C(_10_), .Y(_17_) );
NAND3X1 NAND3X1_683 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_16_), .C(_17_), .Y(_18_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_3767_), .B(bloque_datos[24]), .Y(_19_) );
NAND2X1 NAND2X1_360 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[24]), .B(_3767_), .Y(_20_) );
NAND2X1 NAND2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_19_), .Y(_21_) );
INVX2 INVX2_102 ( .gnd(gnd), .vdd(vdd), .A(_21_), .Y(_22_) );
XNOR2X1 XNOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .B(_22_), .Y(_23_) );
INVX1 INVX1_392 ( .gnd(gnd), .vdd(vdd), .A(_23_), .Y(_24_) );
NAND3X1 NAND3X1_684 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_14_), .C(_18_), .Y(_25_) );
AOI21X1 AOI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_17_), .C(_15_), .Y(_26_) );
AOI21X1 AOI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_9_), .C(_3689_), .Y(_27_) );
OAI21X1 OAI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_27_), .C(_23_), .Y(_28_) );
AOI21X1 AOI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_28_), .C(_3688_), .Y(_29_) );
NAND3X1 NAND3X1_685 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_14_), .C(_18_), .Y(_30_) );
OAI21X1 OAI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_27_), .C(_24_), .Y(_31_) );
AOI21X1 AOI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_31_), .C(bloque_datos[52]), .Y(_32_) );
OAI21X1 OAI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_32_), .C(_3558_), .Y(_33_) );
INVX2 INVX2_103 ( .gnd(gnd), .vdd(vdd), .A(_3558_), .Y(_34_) );
NAND3X1 NAND3X1_686 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[52]), .B(_30_), .C(_31_), .Y(_35_) );
NAND3X1 NAND3X1_687 ( .gnd(gnd), .vdd(vdd), .A(_3688_), .B(_25_), .C(_28_), .Y(_36_) );
NAND3X1 NAND3X1_688 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_35_), .C(_36_), .Y(_37_) );
NAND3X1 NAND3X1_689 ( .gnd(gnd), .vdd(vdd), .A(_3687_), .B(_37_), .C(_33_), .Y(_38_) );
INVX2 INVX2_104 ( .gnd(gnd), .vdd(vdd), .A(_3687_), .Y(_39_) );
NAND3X1 NAND3X1_690 ( .gnd(gnd), .vdd(vdd), .A(_3558_), .B(_35_), .C(_36_), .Y(_40_) );
OAI21X1 OAI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_32_), .C(_34_), .Y(_41_) );
NAND3X1 NAND3X1_691 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_41_), .C(_39_), .Y(_42_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(bloque_datos[40]), .Y(_43_) );
NAND2X1 NAND2X1_362 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[40]), .B(_21_), .Y(_44_) );
NAND2X1 NAND2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_43_), .Y(_45_) );
INVX2 INVX2_105 ( .gnd(gnd), .vdd(vdd), .A(_45_), .Y(_46_) );
XNOR2X1 XNOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1961_), .B(_46_), .Y(_47_) );
INVX1 INVX1_393 ( .gnd(gnd), .vdd(vdd), .A(_47_), .Y(_48_) );
NAND3X1 NAND3X1_692 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_38_), .C(_42_), .Y(_49_) );
AOI21X1 AOI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_41_), .C(_39_), .Y(_50_) );
AOI21X1 AOI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_33_), .C(_3687_), .Y(_51_) );
OAI21X1 OAI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_51_), .C(_47_), .Y(_52_) );
AOI21X1 AOI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_52_), .C(_3686_), .Y(_53_) );
NAND3X1 NAND3X1_693 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_38_), .C(_42_), .Y(_54_) );
OAI21X1 OAI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_51_), .C(_48_), .Y(_55_) );
AOI21X1 AOI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_55_), .C(bloque_datos[68]), .Y(_56_) );
OAI21X1 OAI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_56_), .C(_3574_), .Y(_57_) );
INVX2 INVX2_106 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .Y(_58_) );
NAND3X1 NAND3X1_694 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[68]), .B(_54_), .C(_55_), .Y(_59_) );
NAND3X1 NAND3X1_695 ( .gnd(gnd), .vdd(vdd), .A(_3686_), .B(_49_), .C(_52_), .Y(_60_) );
NAND3X1 NAND3X1_696 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_59_), .C(_60_), .Y(_61_) );
NAND3X1 NAND3X1_697 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_3685_), .C(_57_), .Y(_62_) );
INVX2 INVX2_107 ( .gnd(gnd), .vdd(vdd), .A(_3685_), .Y(_63_) );
NAND3X1 NAND3X1_698 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .B(_59_), .C(_60_), .Y(_64_) );
OAI21X1 OAI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_56_), .C(_58_), .Y(_65_) );
NAND3X1 NAND3X1_699 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_63_), .C(_65_), .Y(_66_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(bloque_datos[56]), .Y(_67_) );
NAND2X1 NAND2X1_364 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[56]), .B(_45_), .Y(_68_) );
NAND2X1 NAND2X1_365 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_67_), .Y(_69_) );
INVX2 INVX2_108 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_70_) );
XNOR2X1 XNOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1994_), .B(_70_), .Y(_71_) );
INVX1 INVX1_394 ( .gnd(gnd), .vdd(vdd), .A(_71_), .Y(_72_) );
NAND3X1 NAND3X1_700 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_66_), .C(_62_), .Y(_73_) );
AOI21X1 AOI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_65_), .C(_63_), .Y(_74_) );
AOI21X1 AOI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_57_), .C(_3685_), .Y(_75_) );
OAI21X1 OAI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_75_), .C(_71_), .Y(_76_) );
AOI21X1 AOI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_76_), .C(_3683_), .Y(_77_) );
NAND3X1 NAND3X1_701 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_66_), .C(_62_), .Y(_78_) );
OAI21X1 OAI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_75_), .C(_72_), .Y(_79_) );
AOI21X1 AOI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_79_), .C(bloque_datos[84]), .Y(_80_) );
OAI21X1 OAI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_80_), .C(_3580_), .Y(_81_) );
INVX2 INVX2_109 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .Y(_82_) );
NAND3X1 NAND3X1_702 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[84]), .B(_78_), .C(_79_), .Y(_83_) );
NAND3X1 NAND3X1_703 ( .gnd(gnd), .vdd(vdd), .A(_3683_), .B(_73_), .C(_76_), .Y(_84_) );
NAND3X1 NAND3X1_704 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_83_), .C(_84_), .Y(_85_) );
NAND3X1 NAND3X1_705 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .B(_85_), .C(_81_), .Y(_86_) );
INVX2 INVX2_110 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .Y(_87_) );
NAND3X1 NAND3X1_706 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_83_), .C(_84_), .Y(_88_) );
OAI21X1 OAI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_80_), .C(_82_), .Y(_89_) );
NAND3X1 NAND3X1_707 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_88_), .C(_89_), .Y(_90_) );
NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[72]), .B(_70_), .Y(_91_) );
NAND2X1 NAND2X1_366 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[72]), .B(_70_), .Y(_92_) );
INVX1 INVX1_395 ( .gnd(gnd), .vdd(vdd), .A(_92_), .Y(_93_) );
NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_93_), .Y(_94_) );
XOR2X1 XOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_2027_), .Y(_95_) );
INVX1 INVX1_396 ( .gnd(gnd), .vdd(vdd), .A(_95_), .Y(_96_) );
NAND3X1 NAND3X1_708 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_86_), .C(_90_), .Y(_97_) );
AOI21X1 AOI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_89_), .C(_87_), .Y(_98_) );
AOI21X1 AOI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_81_), .C(_3682_), .Y(_99_) );
OAI21X1 OAI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_99_), .C(_95_), .Y(_100_) );
AOI21X1 AOI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_100_), .C(_3681_), .Y(_101_) );
NAND3X1 NAND3X1_709 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_86_), .C(_90_), .Y(_102_) );
OAI21X1 OAI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_99_), .C(_96_), .Y(_103_) );
AOI21X1 AOI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_103_), .C(W_132_), .Y(_104_) );
OAI21X1 OAI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_104_), .C(_3595_), .Y(_105_) );
INVX2 INVX2_111 ( .gnd(gnd), .vdd(vdd), .A(_3595_), .Y(_106_) );
NAND3X1 NAND3X1_710 ( .gnd(gnd), .vdd(vdd), .A(W_132_), .B(_102_), .C(_103_), .Y(_107_) );
NAND3X1 NAND3X1_711 ( .gnd(gnd), .vdd(vdd), .A(_3681_), .B(_97_), .C(_100_), .Y(_108_) );
NAND3X1 NAND3X1_712 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_107_), .C(_108_), .Y(_109_) );
NAND3X1 NAND3X1_713 ( .gnd(gnd), .vdd(vdd), .A(_3680_), .B(_109_), .C(_105_), .Y(_110_) );
NAND3X1 NAND3X1_714 ( .gnd(gnd), .vdd(vdd), .A(_3595_), .B(_107_), .C(_108_), .Y(_111_) );
OAI21X1 OAI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_104_), .C(_106_), .Y(_112_) );
NAND3X1 NAND3X1_715 ( .gnd(gnd), .vdd(vdd), .A(_3679_), .B(_111_), .C(_112_), .Y(_113_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(bloque_datos[88]), .Y(_114_) );
NAND2X1 NAND2X1_367 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .B(_94_), .Y(_115_) );
NAND2X1 NAND2X1_368 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_114_), .Y(_116_) );
NAND3X1 NAND3X1_716 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_110_), .C(_113_), .Y(_117_) );
AOI21X1 AOI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_112_), .C(_3679_), .Y(_118_) );
AOI21X1 AOI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_105_), .C(_3680_), .Y(_119_) );
INVX2 INVX2_112 ( .gnd(gnd), .vdd(vdd), .A(_116_), .Y(_120_) );
OAI21X1 OAI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_119_), .C(_120_), .Y(_121_) );
NAND3X1 NAND3X1_717 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(_117_), .C(_121_), .Y(_122_) );
NAND2X1 NAND2X1_369 ( .gnd(gnd), .vdd(vdd), .A(W_148_), .B(_122_), .Y(_123_) );
INVX1 INVX1_397 ( .gnd(gnd), .vdd(vdd), .A(W_148_), .Y(_124_) );
NAND2X1 NAND2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_113_), .Y(_125_) );
AOI21X1 AOI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_125_), .C(_2411_), .Y(_126_) );
NAND3X1 NAND3X1_718 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_117_), .C(_126_), .Y(_127_) );
NAND3X1 NAND3X1_719 ( .gnd(gnd), .vdd(vdd), .A(_3678_), .B(_127_), .C(_123_), .Y(_128_) );
NAND2X1 NAND2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_122_), .Y(_129_) );
NAND3X1 NAND3X1_720 ( .gnd(gnd), .vdd(vdd), .A(W_148_), .B(_117_), .C(_126_), .Y(_130_) );
NAND3X1 NAND3X1_721 ( .gnd(gnd), .vdd(vdd), .A(_3604_), .B(_130_), .C(_129_), .Y(_131_) );
NAND3X1 NAND3X1_722 ( .gnd(gnd), .vdd(vdd), .A(_3677_), .B(_128_), .C(_131_), .Y(_132_) );
INVX2 INVX2_113 ( .gnd(gnd), .vdd(vdd), .A(_3677_), .Y(_133_) );
AOI21X1 AOI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_129_), .C(_3604_), .Y(_134_) );
AOI21X1 AOI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_123_), .C(_3678_), .Y(_135_) );
OAI21X1 OAI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_135_), .C(_133_), .Y(_136_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(W_136_), .Y(_137_) );
NAND2X1 NAND2X1_372 ( .gnd(gnd), .vdd(vdd), .A(W_136_), .B(_116_), .Y(_138_) );
NAND2X1 NAND2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_137_), .Y(_139_) );
NAND3X1 NAND3X1_723 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_139_), .C(_136_), .Y(_140_) );
NOR3X1 NOR3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_133_), .C(_135_), .Y(_141_) );
AOI21X1 AOI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_131_), .C(_3677_), .Y(_142_) );
INVX2 INVX2_114 ( .gnd(gnd), .vdd(vdd), .A(_139_), .Y(_143_) );
OAI21X1 OAI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_142_), .C(_143_), .Y(_144_) );
NAND3X1 NAND3X1_724 ( .gnd(gnd), .vdd(vdd), .A(_2093_), .B(_140_), .C(_144_), .Y(_145_) );
NAND2X1 NAND2X1_374 ( .gnd(gnd), .vdd(vdd), .A(W_164_), .B(_145_), .Y(_146_) );
INVX1 INVX1_398 ( .gnd(gnd), .vdd(vdd), .A(W_164_), .Y(_147_) );
OAI21X1 OAI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_142_), .C(_139_), .Y(_148_) );
NAND3X1 NAND3X1_725 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_143_), .C(_136_), .Y(_149_) );
NAND2X1 NAND2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_148_), .Y(_150_) );
NAND3X1 NAND3X1_726 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_2093_), .C(_150_), .Y(_151_) );
NAND3X1 NAND3X1_727 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .B(_146_), .C(_151_), .Y(_152_) );
NAND2X1 NAND2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_145_), .Y(_153_) );
NAND3X1 NAND3X1_728 ( .gnd(gnd), .vdd(vdd), .A(W_164_), .B(_2093_), .C(_150_), .Y(_154_) );
NAND3X1 NAND3X1_729 ( .gnd(gnd), .vdd(vdd), .A(_3674_), .B(_153_), .C(_154_), .Y(_155_) );
NAND3X1 NAND3X1_730 ( .gnd(gnd), .vdd(vdd), .A(_3672_), .B(_152_), .C(_155_), .Y(_156_) );
INVX2 INVX2_115 ( .gnd(gnd), .vdd(vdd), .A(_3672_), .Y(_157_) );
AOI21X1 AOI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_154_), .C(_3674_), .Y(_158_) );
AOI21X1 AOI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_151_), .C(_3675_), .Y(_159_) );
OAI21X1 OAI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_159_), .C(_157_), .Y(_160_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(W_152_), .Y(_161_) );
NAND2X1 NAND2X1_377 ( .gnd(gnd), .vdd(vdd), .A(W_152_), .B(_139_), .Y(_162_) );
NAND2X1 NAND2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_161_), .Y(_163_) );
NAND3X1 NAND3X1_731 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_163_), .C(_160_), .Y(_164_) );
NOR3X1 NOR3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_157_), .C(_159_), .Y(_165_) );
AOI21X1 AOI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_155_), .C(_3672_), .Y(_166_) );
INVX2 INVX2_116 ( .gnd(gnd), .vdd(vdd), .A(_163_), .Y(_167_) );
OAI21X1 OAI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_166_), .C(_167_), .Y(_168_) );
NAND3X1 NAND3X1_732 ( .gnd(gnd), .vdd(vdd), .A(_2126_), .B(_164_), .C(_168_), .Y(_169_) );
NAND2X1 NAND2X1_379 ( .gnd(gnd), .vdd(vdd), .A(W_180_), .B(_169_), .Y(_170_) );
INVX1 INVX1_399 ( .gnd(gnd), .vdd(vdd), .A(W_180_), .Y(_171_) );
OAI21X1 OAI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_166_), .C(_163_), .Y(_172_) );
NAND3X1 NAND3X1_733 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_167_), .C(_160_), .Y(_173_) );
NAND2X1 NAND2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_172_), .Y(_174_) );
NAND3X1 NAND3X1_734 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_2126_), .C(_174_), .Y(_175_) );
NAND3X1 NAND3X1_735 ( .gnd(gnd), .vdd(vdd), .A(_3671_), .B(_170_), .C(_175_), .Y(_176_) );
NAND2X1 NAND2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_169_), .Y(_177_) );
NAND3X1 NAND3X1_736 ( .gnd(gnd), .vdd(vdd), .A(W_180_), .B(_2126_), .C(_174_), .Y(_178_) );
NAND3X1 NAND3X1_737 ( .gnd(gnd), .vdd(vdd), .A(_3670_), .B(_177_), .C(_178_), .Y(_179_) );
NAND3X1 NAND3X1_738 ( .gnd(gnd), .vdd(vdd), .A(_3668_), .B(_176_), .C(_179_), .Y(_180_) );
INVX2 INVX2_117 ( .gnd(gnd), .vdd(vdd), .A(_3668_), .Y(_181_) );
AOI21X1 AOI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_178_), .C(_3670_), .Y(_182_) );
AOI21X1 AOI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_175_), .C(_3671_), .Y(_183_) );
OAI21X1 OAI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_183_), .C(_181_), .Y(_184_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(W_168_), .Y(_185_) );
NAND2X1 NAND2X1_382 ( .gnd(gnd), .vdd(vdd), .A(W_168_), .B(_163_), .Y(_186_) );
NAND2X1 NAND2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_185_), .Y(_187_) );
NAND3X1 NAND3X1_739 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_187_), .C(_184_), .Y(_188_) );
NOR3X1 NOR3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_181_), .C(_183_), .Y(_189_) );
AOI21X1 AOI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_179_), .C(_3668_), .Y(_190_) );
INVX2 INVX2_118 ( .gnd(gnd), .vdd(vdd), .A(_187_), .Y(_191_) );
OAI21X1 OAI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_190_), .C(_191_), .Y(_192_) );
NAND3X1 NAND3X1_740 ( .gnd(gnd), .vdd(vdd), .A(_2159_), .B(_188_), .C(_192_), .Y(_193_) );
NAND2X1 NAND2X1_384 ( .gnd(gnd), .vdd(vdd), .A(W_196_), .B(_193_), .Y(_194_) );
INVX1 INVX1_400 ( .gnd(gnd), .vdd(vdd), .A(W_196_), .Y(_195_) );
OAI21X1 OAI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_190_), .C(_187_), .Y(_196_) );
NAND3X1 NAND3X1_741 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_191_), .C(_184_), .Y(_197_) );
NAND2X1 NAND2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_196_), .Y(_198_) );
NAND3X1 NAND3X1_742 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_2159_), .C(_198_), .Y(_199_) );
NAND3X1 NAND3X1_743 ( .gnd(gnd), .vdd(vdd), .A(_3666_), .B(_194_), .C(_199_), .Y(_200_) );
NAND2X1 NAND2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_193_), .Y(_201_) );
NAND3X1 NAND3X1_744 ( .gnd(gnd), .vdd(vdd), .A(W_196_), .B(_2159_), .C(_198_), .Y(_202_) );
NAND3X1 NAND3X1_745 ( .gnd(gnd), .vdd(vdd), .A(_3665_), .B(_201_), .C(_202_), .Y(_203_) );
NAND3X1 NAND3X1_746 ( .gnd(gnd), .vdd(vdd), .A(_3663_), .B(_200_), .C(_203_), .Y(_204_) );
INVX2 INVX2_119 ( .gnd(gnd), .vdd(vdd), .A(_3663_), .Y(_205_) );
AOI21X1 AOI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_202_), .C(_3665_), .Y(_206_) );
AOI21X1 AOI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_199_), .C(_3666_), .Y(_207_) );
OAI21X1 OAI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_207_), .C(_205_), .Y(_208_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(W_184_), .Y(_209_) );
NAND2X1 NAND2X1_387 ( .gnd(gnd), .vdd(vdd), .A(W_184_), .B(_187_), .Y(_210_) );
NAND2X1 NAND2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_210_), .B(_209_), .Y(_211_) );
NAND3X1 NAND3X1_747 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_211_), .C(_208_), .Y(_212_) );
NAND3X1 NAND3X1_748 ( .gnd(gnd), .vdd(vdd), .A(_3665_), .B(_194_), .C(_199_), .Y(_213_) );
NAND3X1 NAND3X1_749 ( .gnd(gnd), .vdd(vdd), .A(_3666_), .B(_201_), .C(_202_), .Y(_214_) );
AOI21X1 AOI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_214_), .C(_205_), .Y(_215_) );
AOI21X1 AOI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_203_), .C(_3663_), .Y(_216_) );
INVX2 INVX2_120 ( .gnd(gnd), .vdd(vdd), .A(_211_), .Y(_217_) );
OAI21X1 OAI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_216_), .C(_217_), .Y(_218_) );
NAND3X1 NAND3X1_750 ( .gnd(gnd), .vdd(vdd), .A(_2192_), .B(_212_), .C(_218_), .Y(_219_) );
NAND2X1 NAND2X1_389 ( .gnd(gnd), .vdd(vdd), .A(W_212_), .B(_219_), .Y(_220_) );
INVX1 INVX1_401 ( .gnd(gnd), .vdd(vdd), .A(W_212_), .Y(_221_) );
OAI21X1 OAI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_216_), .C(_211_), .Y(_222_) );
NAND3X1 NAND3X1_751 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_217_), .C(_208_), .Y(_223_) );
NAND2X1 NAND2X1_390 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_222_), .Y(_224_) );
NAND3X1 NAND3X1_752 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_2192_), .C(_224_), .Y(_225_) );
NAND3X1 NAND3X1_753 ( .gnd(gnd), .vdd(vdd), .A(_3662_), .B(_220_), .C(_225_), .Y(_226_) );
NAND2X1 NAND2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_219_), .Y(_227_) );
NAND3X1 NAND3X1_754 ( .gnd(gnd), .vdd(vdd), .A(W_212_), .B(_2192_), .C(_224_), .Y(_228_) );
NAND3X1 NAND3X1_755 ( .gnd(gnd), .vdd(vdd), .A(_3661_), .B(_227_), .C(_228_), .Y(_229_) );
NAND3X1 NAND3X1_756 ( .gnd(gnd), .vdd(vdd), .A(_3659_), .B(_226_), .C(_229_), .Y(_230_) );
AOI21X1 AOI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_228_), .C(_3661_), .Y(_231_) );
AOI21X1 AOI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_225_), .C(_3662_), .Y(_232_) );
OAI21X1 OAI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_232_), .C(_3658_), .Y(_233_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(W_200_), .Y(_234_) );
NAND2X1 NAND2X1_392 ( .gnd(gnd), .vdd(vdd), .A(W_200_), .B(_211_), .Y(_235_) );
NAND2X1 NAND2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_234_), .Y(_236_) );
NAND3X1 NAND3X1_757 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_236_), .C(_233_), .Y(_237_) );
NAND3X1 NAND3X1_758 ( .gnd(gnd), .vdd(vdd), .A(_3661_), .B(_220_), .C(_225_), .Y(_238_) );
NAND3X1 NAND3X1_759 ( .gnd(gnd), .vdd(vdd), .A(_3662_), .B(_227_), .C(_228_), .Y(_239_) );
AOI21X1 AOI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_239_), .C(_3658_), .Y(_240_) );
AOI21X1 AOI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_229_), .C(_3659_), .Y(_241_) );
INVX2 INVX2_121 ( .gnd(gnd), .vdd(vdd), .A(_236_), .Y(_242_) );
OAI21X1 OAI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_241_), .C(_242_), .Y(_243_) );
NAND3X1 NAND3X1_760 ( .gnd(gnd), .vdd(vdd), .A(_2225_), .B(_237_), .C(_243_), .Y(_244_) );
NAND2X1 NAND2X1_394 ( .gnd(gnd), .vdd(vdd), .A(W_228_), .B(_244_), .Y(_245_) );
INVX1 INVX1_402 ( .gnd(gnd), .vdd(vdd), .A(W_228_), .Y(_246_) );
OAI21X1 OAI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_241_), .C(_236_), .Y(_247_) );
NAND3X1 NAND3X1_761 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_242_), .C(_233_), .Y(_248_) );
AOI21X1 AOI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_247_), .C(_2290_), .Y(_249_) );
NAND2X1 NAND2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_249_), .Y(_250_) );
NAND3X1 NAND3X1_762 ( .gnd(gnd), .vdd(vdd), .A(_3656_), .B(_245_), .C(_250_), .Y(_251_) );
NAND2X1 NAND2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_244_), .Y(_252_) );
NAND2X1 NAND2X1_397 ( .gnd(gnd), .vdd(vdd), .A(W_228_), .B(_249_), .Y(_253_) );
NAND3X1 NAND3X1_763 ( .gnd(gnd), .vdd(vdd), .A(_3655_), .B(_252_), .C(_253_), .Y(_254_) );
NAND3X1 NAND3X1_764 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_254_), .C(_3653_), .Y(_255_) );
AOI21X1 AOI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_253_), .C(_3655_), .Y(_256_) );
AOI21X1 AOI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_250_), .C(_3656_), .Y(_257_) );
OAI21X1 OAI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_257_), .C(_3652_), .Y(_258_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(W_216_), .Y(_259_) );
NAND2X1 NAND2X1_398 ( .gnd(gnd), .vdd(vdd), .A(W_216_), .B(_236_), .Y(_260_) );
NAND2X1 NAND2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_259_), .Y(_261_) );
NAND3X1 NAND3X1_765 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_255_), .C(_258_), .Y(_262_) );
NOR3X1 NOR3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_3652_), .C(_257_), .Y(_263_) );
AOI21X1 AOI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_254_), .C(_3653_), .Y(_264_) );
INVX2 INVX2_122 ( .gnd(gnd), .vdd(vdd), .A(_261_), .Y(_265_) );
OAI21X1 OAI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_264_), .C(_265_), .Y(_266_) );
NAND3X1 NAND3X1_766 ( .gnd(gnd), .vdd(vdd), .A(_2257_), .B(_262_), .C(_266_), .Y(_267_) );
NAND2X1 NAND2X1_400 ( .gnd(gnd), .vdd(vdd), .A(W_244_), .B(_267_), .Y(_268_) );
INVX1 INVX1_403 ( .gnd(gnd), .vdd(vdd), .A(W_244_), .Y(_269_) );
NAND2X1 NAND2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_258_), .Y(_270_) );
AOI21X1 AOI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_270_), .C(_2268_), .Y(_271_) );
NAND3X1 NAND3X1_767 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_262_), .C(_271_), .Y(_272_) );
NAND3X1 NAND3X1_768 ( .gnd(gnd), .vdd(vdd), .A(_3642_), .B(_272_), .C(_268_), .Y(_273_) );
INVX1 INVX1_404 ( .gnd(gnd), .vdd(vdd), .A(_3642_), .Y(_274_) );
NAND2X1 NAND2X1_402 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_267_), .Y(_275_) );
NAND3X1 NAND3X1_769 ( .gnd(gnd), .vdd(vdd), .A(W_244_), .B(_262_), .C(_271_), .Y(_276_) );
NAND3X1 NAND3X1_770 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_276_), .C(_275_), .Y(_277_) );
NAND3X1 NAND3X1_771 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_277_), .C(_3651_), .Y(_278_) );
INVX1 INVX1_405 ( .gnd(gnd), .vdd(vdd), .A(_3646_), .Y(_279_) );
AOI21X1 AOI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3472_), .C(_279_), .Y(_280_) );
AOI21X1 AOI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_275_), .C(_274_), .Y(_281_) );
AOI21X1 AOI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_268_), .C(_3642_), .Y(_282_) );
OAI21X1 OAI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_282_), .C(_280_), .Y(_283_) );
NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(W_232_), .B(_265_), .Y(_284_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(W_232_), .Y(_285_) );
NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_285_), .Y(_286_) );
INVX2 INVX2_123 ( .gnd(gnd), .vdd(vdd), .A(_286_), .Y(_287_) );
NAND3X1 NAND3X1_772 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_287_), .C(_278_), .Y(_288_) );
NOR3X1 NOR3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_282_), .C(_280_), .Y(_289_) );
AOI21X1 AOI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_277_), .C(_3651_), .Y(_290_) );
OAI21X1 OAI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_290_), .C(_286_), .Y(_291_) );
NAND3X1 NAND3X1_773 ( .gnd(gnd), .vdd(vdd), .A(_3648_), .B(_288_), .C(_291_), .Y(_292_) );
INVX1 INVX1_406 ( .gnd(gnd), .vdd(vdd), .A(_292_), .Y(_293_) );
AOI21X1 AOI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_291_), .C(_3648_), .Y(_294_) );
NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_293_), .Y(H_4_) );
INVX1 INVX1_407 ( .gnd(gnd), .vdd(vdd), .A(W_233_), .Y(_295_) );
INVX1 INVX1_408 ( .gnd(gnd), .vdd(vdd), .A(W_217_), .Y(_296_) );
INVX1 INVX1_409 ( .gnd(gnd), .vdd(vdd), .A(W_201_), .Y(_297_) );
INVX1 INVX1_410 ( .gnd(gnd), .vdd(vdd), .A(W_185_), .Y(_298_) );
INVX1 INVX1_411 ( .gnd(gnd), .vdd(vdd), .A(W_169_), .Y(_299_) );
INVX1 INVX1_412 ( .gnd(gnd), .vdd(vdd), .A(W_153_), .Y(_300_) );
NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(W_136_), .B(_120_), .Y(_301_) );
INVX1 INVX1_413 ( .gnd(gnd), .vdd(vdd), .A(_94_), .Y(_302_) );
NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .B(_302_), .Y(_303_) );
NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[56]), .B(_46_), .Y(_304_) );
INVX1 INVX1_414 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[57]), .Y(_305_) );
NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[40]), .B(_22_), .Y(_306_) );
INVX1 INVX1_415 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[41]), .Y(_307_) );
NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[24]), .B(_3768_), .Y(_308_) );
INVX1 INVX1_416 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[25]), .Y(_309_) );
NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .B(_3742_), .Y(_310_) );
INVX1 INVX1_417 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .Y(_311_) );
NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(W_25_), .B(W_9_), .Y(_312_) );
INVX1 INVX1_418 ( .gnd(gnd), .vdd(vdd), .A(W_25_), .Y(_313_) );
INVX2 INVX2_124 ( .gnd(gnd), .vdd(vdd), .A(W_9_), .Y(_314_) );
NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_314_), .Y(_315_) );
NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_315_), .Y(_316_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_3740_), .Y(_317_) );
NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_3740_), .B(_316_), .Y(_318_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_318_), .Y(_319_) );
NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_319_), .Y(_320_) );
NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_317_), .Y(_321_) );
NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .B(_321_), .Y(_322_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_322_), .Y(_323_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_310_), .Y(_324_) );
OAI21X1 OAI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_322_), .C(_310_), .Y(_325_) );
NAND2X1 NAND2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_324_), .Y(_326_) );
NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_326_), .Y(_327_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_325_), .Y(_328_) );
NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[25]), .B(_328_), .Y(_329_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_327_), .Y(_330_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_308_), .Y(_331_) );
OAI21X1 OAI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_327_), .C(_308_), .Y(_332_) );
NAND2X1 NAND2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_331_), .Y(_333_) );
NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_333_), .Y(_334_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_332_), .Y(_335_) );
NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[41]), .B(_335_), .Y(_336_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_334_), .Y(_337_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_306_), .Y(_338_) );
OAI21X1 OAI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_334_), .C(_306_), .Y(_339_) );
NAND2X1 NAND2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_338_), .Y(_340_) );
NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_340_), .Y(_341_) );
AOI21X1 AOI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_338_), .C(bloque_datos[57]), .Y(_342_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_342_), .Y(_343_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_304_), .Y(_344_) );
OAI21X1 OAI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_342_), .C(_304_), .Y(_345_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_345_), .Y(_346_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(bloque_datos[73]), .Y(_347_) );
NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[73]), .B(_346_), .Y(_348_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_348_), .Y(_349_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_91_), .Y(_350_) );
OAI21X1 OAI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_348_), .C(_91_), .Y(_351_) );
NAND2X1 NAND2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_350_), .Y(_352_) );
INVX2 INVX2_125 ( .gnd(gnd), .vdd(vdd), .A(_352_), .Y(_353_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(bloque_datos[89]), .Y(_354_) );
NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[89]), .B(_353_), .Y(_355_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_355_), .Y(_356_) );
NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_356_), .Y(_357_) );
INVX2 INVX2_126 ( .gnd(gnd), .vdd(vdd), .A(_357_), .Y(_358_) );
OAI21X1 OAI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_355_), .C(_303_), .Y(_359_) );
NAND2X1 NAND2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_358_), .Y(_360_) );
INVX2 INVX2_127 ( .gnd(gnd), .vdd(vdd), .A(_360_), .Y(_361_) );
NAND2X1 NAND2X1_408 ( .gnd(gnd), .vdd(vdd), .A(W_137_), .B(_361_), .Y(_362_) );
INVX1 INVX1_419 ( .gnd(gnd), .vdd(vdd), .A(W_137_), .Y(_363_) );
NAND2X1 NAND2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_360_), .Y(_364_) );
NAND2X1 NAND2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_362_), .Y(_365_) );
NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_365_), .Y(_366_) );
INVX1 INVX1_420 ( .gnd(gnd), .vdd(vdd), .A(_366_), .Y(_367_) );
NAND2X1 NAND2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_365_), .Y(_368_) );
NAND2X1 NAND2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_367_), .Y(_369_) );
NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_369_), .Y(_370_) );
INVX2 INVX2_128 ( .gnd(gnd), .vdd(vdd), .A(_370_), .Y(_371_) );
NAND2X1 NAND2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_369_), .Y(_372_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_372_), .Y(_373_) );
OAI21X1 OAI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(W_152_), .B(_143_), .C(_373_), .Y(_374_) );
NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(W_152_), .B(_143_), .Y(_375_) );
INVX1 INVX1_421 ( .gnd(gnd), .vdd(vdd), .A(_373_), .Y(_376_) );
NAND2X1 NAND2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_376_), .Y(_377_) );
NAND2X1 NAND2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_377_), .Y(_378_) );
NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_378_), .Y(_379_) );
INVX2 INVX2_129 ( .gnd(gnd), .vdd(vdd), .A(_378_), .Y(_380_) );
NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(W_169_), .B(_380_), .Y(_381_) );
NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_381_), .Y(_382_) );
OAI21X1 OAI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(W_168_), .B(_167_), .C(_382_), .Y(_383_) );
NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(W_168_), .B(_167_), .Y(_384_) );
OAI21X1 OAI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_379_), .C(_384_), .Y(_385_) );
NAND2X1 NAND2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_383_), .Y(_386_) );
NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_386_), .Y(_387_) );
INVX2 INVX2_130 ( .gnd(gnd), .vdd(vdd), .A(_386_), .Y(_388_) );
NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(W_185_), .B(_388_), .Y(_389_) );
NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_389_), .Y(_390_) );
OAI21X1 OAI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(W_184_), .B(_191_), .C(_390_), .Y(_391_) );
NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(W_184_), .B(_191_), .Y(_392_) );
OAI21X1 OAI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_387_), .C(_392_), .Y(_393_) );
NAND2X1 NAND2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_391_), .Y(_394_) );
NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_394_), .Y(_395_) );
INVX2 INVX2_131 ( .gnd(gnd), .vdd(vdd), .A(_394_), .Y(_396_) );
NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(W_201_), .B(_396_), .Y(_397_) );
NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_397_), .Y(_398_) );
OAI21X1 OAI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(W_200_), .B(_217_), .C(_398_), .Y(_399_) );
NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(W_200_), .B(_217_), .Y(_400_) );
OAI21X1 OAI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_395_), .C(_400_), .Y(_401_) );
NAND2X1 NAND2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_399_), .Y(_402_) );
NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_402_), .Y(_403_) );
INVX2 INVX2_132 ( .gnd(gnd), .vdd(vdd), .A(_402_), .Y(_404_) );
NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(W_217_), .B(_404_), .Y(_405_) );
NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_405_), .Y(_406_) );
OAI21X1 OAI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(W_216_), .B(_242_), .C(_406_), .Y(_407_) );
NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(W_216_), .B(_242_), .Y(_408_) );
OAI21X1 OAI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_403_), .C(_408_), .Y(_409_) );
NAND2X1 NAND2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_407_), .Y(_410_) );
NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_410_), .Y(_411_) );
INVX1 INVX1_422 ( .gnd(gnd), .vdd(vdd), .A(_410_), .Y(_412_) );
NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(W_233_), .B(_412_), .Y(_413_) );
NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_413_), .Y(_414_) );
OAI21X1 OAI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(W_232_), .B(_265_), .C(_414_), .Y(_415_) );
OAI21X1 OAI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_411_), .C(_284_), .Y(_416_) );
NAND2X1 NAND2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_415_), .Y(_417_) );
INVX2 INVX2_133 ( .gnd(gnd), .vdd(vdd), .A(_417_), .Y(_418_) );
OAI21X1 OAI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_282_), .C(_273_), .Y(_419_) );
OAI21X1 OAI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_3652_), .C(_251_), .Y(_420_) );
INVX2 INVX2_134 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_421_) );
INVX1 INVX1_423 ( .gnd(gnd), .vdd(vdd), .A(W_229_), .Y(_422_) );
OAI21X1 OAI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_3658_), .C(_226_), .Y(_423_) );
INVX2 INVX2_135 ( .gnd(gnd), .vdd(vdd), .A(_220_), .Y(_424_) );
INVX1 INVX1_424 ( .gnd(gnd), .vdd(vdd), .A(W_213_), .Y(_425_) );
OAI21X1 OAI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_205_), .C(_200_), .Y(_426_) );
INVX2 INVX2_136 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(_427_) );
INVX1 INVX1_425 ( .gnd(gnd), .vdd(vdd), .A(W_197_), .Y(_428_) );
OAI21X1 OAI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_181_), .C(_176_), .Y(_429_) );
INVX1 INVX1_426 ( .gnd(gnd), .vdd(vdd), .A(_170_), .Y(_430_) );
INVX1 INVX1_427 ( .gnd(gnd), .vdd(vdd), .A(W_181_), .Y(_431_) );
OAI21X1 OAI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(_157_), .C(_152_), .Y(_432_) );
INVX1 INVX1_428 ( .gnd(gnd), .vdd(vdd), .A(_146_), .Y(_433_) );
INVX1 INVX1_429 ( .gnd(gnd), .vdd(vdd), .A(W_165_), .Y(_434_) );
OAI21X1 OAI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_133_), .C(_128_), .Y(_435_) );
INVX1 INVX1_430 ( .gnd(gnd), .vdd(vdd), .A(_123_), .Y(_436_) );
INVX1 INVX1_431 ( .gnd(gnd), .vdd(vdd), .A(W_149_), .Y(_437_) );
NOR3X1 NOR3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_3595_), .C(_104_), .Y(_438_) );
OAI21X1 OAI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_3679_), .C(_105_), .Y(_439_) );
NOR3X1 NOR3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_3580_), .C(_80_), .Y(_440_) );
OAI21X1 OAI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_87_), .C(_81_), .Y(_441_) );
NOR3X1 NOR3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_3574_), .C(_56_), .Y(_442_) );
OAI21X1 OAI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_63_), .C(_57_), .Y(_443_) );
NOR3X1 NOR3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_3558_), .C(_32_), .Y(_444_) );
OAI21X1 OAI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_39_), .C(_33_), .Y(_445_) );
NAND2X1 NAND2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_14_), .Y(_446_) );
NAND2X1 NAND2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_3753_), .B(_3758_), .Y(_447_) );
INVX1 INVX1_432 ( .gnd(gnd), .vdd(vdd), .A(_3736_), .Y(_448_) );
AOI21X1 AOI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_3737_), .B(_3735_), .C(_448_), .Y(_449_) );
INVX1 INVX1_433 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[5]), .Y(_450_) );
AOI21X1 AOI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_3708_), .B(_3705_), .C(_3508_), .Y(_451_) );
INVX1 INVX1_434 ( .gnd(gnd), .vdd(vdd), .A(W_21_), .Y(_452_) );
NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_2630_), .B(_2674_), .Y(_453_) );
INVX2 INVX2_137 ( .gnd(gnd), .vdd(vdd), .A(W_5_), .Y(_454_) );
XNOR2X1 XNOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(_454_), .Y(_455_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_453_), .Y(_456_) );
NAND2X1 NAND2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_455_), .Y(_457_) );
NAND3X1 NAND3X1_774 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_457_), .C(_456_), .Y(_458_) );
NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(W_5_), .B(_3699_), .Y(_459_) );
NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_3703_), .Y(_460_) );
OAI21X1 OAI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_459_), .C(_453_), .Y(_461_) );
OAI21X1 OAI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_2630_), .B(_2674_), .C(_455_), .Y(_462_) );
NAND3X1 NAND3X1_775 ( .gnd(gnd), .vdd(vdd), .A(W_21_), .B(_462_), .C(_461_), .Y(_463_) );
NAND3X1 NAND3X1_776 ( .gnd(gnd), .vdd(vdd), .A(_3705_), .B(_463_), .C(_458_), .Y(_464_) );
INVX1 INVX1_435 ( .gnd(gnd), .vdd(vdd), .A(_3705_), .Y(_465_) );
NAND3X1 NAND3X1_777 ( .gnd(gnd), .vdd(vdd), .A(W_21_), .B(_457_), .C(_456_), .Y(_466_) );
NAND3X1 NAND3X1_778 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_462_), .C(_461_), .Y(_467_) );
NAND3X1 NAND3X1_779 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_467_), .C(_466_), .Y(_468_) );
NAND2X1 NAND2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_468_), .Y(_469_) );
OAI21X1 OAI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_3723_), .C(_469_), .Y(_470_) );
NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_3723_), .Y(_471_) );
NAND3X1 NAND3X1_780 ( .gnd(gnd), .vdd(vdd), .A(_3705_), .B(_467_), .C(_466_), .Y(_472_) );
NAND3X1 NAND3X1_781 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_463_), .C(_458_), .Y(_473_) );
NAND2X1 NAND2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_473_), .Y(_474_) );
NAND2X1 NAND2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_471_), .Y(_475_) );
XNOR2X1 XNOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_2751_), .B(W_9_), .Y(_476_) );
NAND3X1 NAND3X1_782 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_470_), .C(_475_), .Y(_477_) );
NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_471_), .Y(_478_) );
NAND2X1 NAND2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(_3718_), .Y(_479_) );
NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_479_), .Y(_480_) );
INVX1 INVX1_436 ( .gnd(gnd), .vdd(vdd), .A(_476_), .Y(_481_) );
OAI21X1 OAI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_480_), .C(_481_), .Y(_482_) );
NAND3X1 NAND3X1_783 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_477_), .C(_482_), .Y(_483_) );
NAND3X1 NAND3X1_784 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_470_), .C(_475_), .Y(_484_) );
OAI21X1 OAI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_480_), .C(_476_), .Y(_485_) );
NAND3X1 NAND3X1_785 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[5]), .B(_484_), .C(_485_), .Y(_486_) );
NAND3X1 NAND3X1_786 ( .gnd(gnd), .vdd(vdd), .A(_3729_), .B(_483_), .C(_486_), .Y(_487_) );
NAND3X1 NAND3X1_787 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[5]), .B(_477_), .C(_482_), .Y(_488_) );
NAND3X1 NAND3X1_788 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_484_), .C(_485_), .Y(_489_) );
NAND3X1 NAND3X1_789 ( .gnd(gnd), .vdd(vdd), .A(_3732_), .B(_488_), .C(_489_), .Y(_490_) );
AOI21X1 AOI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_490_), .C(_449_), .Y(_491_) );
NAND2X1 NAND2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_3736_), .B(_3745_), .Y(_492_) );
NAND3X1 NAND3X1_790 ( .gnd(gnd), .vdd(vdd), .A(_3729_), .B(_488_), .C(_489_), .Y(_493_) );
NAND3X1 NAND3X1_791 ( .gnd(gnd), .vdd(vdd), .A(_3732_), .B(_483_), .C(_486_), .Y(_494_) );
AOI21X1 AOI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_494_), .C(_492_), .Y(_495_) );
NAND2X1 NAND2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_2828_), .B(_2795_), .Y(_496_) );
XNOR2X1 XNOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_321_), .Y(_497_) );
NOR3X1 NOR3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_497_), .C(_495_), .Y(_498_) );
NAND3X1 NAND3X1_792 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_494_), .C(_492_), .Y(_499_) );
NAND3X1 NAND3X1_793 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_487_), .C(_490_), .Y(_500_) );
INVX1 INVX1_437 ( .gnd(gnd), .vdd(vdd), .A(_497_), .Y(_501_) );
AOI21X1 AOI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_499_), .C(_501_), .Y(_502_) );
OAI21X1 OAI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_502_), .C(bloque_datos[21]), .Y(_503_) );
INVX1 INVX1_438 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[21]), .Y(_504_) );
NAND3X1 NAND3X1_794 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_500_), .C(_499_), .Y(_505_) );
OAI21X1 OAI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_495_), .C(_497_), .Y(_506_) );
NAND3X1 NAND3X1_795 ( .gnd(gnd), .vdd(vdd), .A(_504_), .B(_505_), .C(_506_), .Y(_507_) );
NAND3X1 NAND3X1_796 ( .gnd(gnd), .vdd(vdd), .A(_3756_), .B(_507_), .C(_503_), .Y(_508_) );
OAI21X1 OAI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_502_), .C(_504_), .Y(_509_) );
NAND3X1 NAND3X1_797 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[21]), .B(_505_), .C(_506_), .Y(_510_) );
NAND3X1 NAND3X1_798 ( .gnd(gnd), .vdd(vdd), .A(_3752_), .B(_510_), .C(_509_), .Y(_511_) );
NAND3X1 NAND3X1_799 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_447_), .C(_511_), .Y(_512_) );
INVX1 INVX1_439 ( .gnd(gnd), .vdd(vdd), .A(_3753_), .Y(_513_) );
AOI21X1 AOI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_3757_), .B(_3692_), .C(_513_), .Y(_514_) );
NAND3X1 NAND3X1_800 ( .gnd(gnd), .vdd(vdd), .A(_3756_), .B(_510_), .C(_509_), .Y(_515_) );
NAND3X1 NAND3X1_801 ( .gnd(gnd), .vdd(vdd), .A(_3752_), .B(_507_), .C(_503_), .Y(_516_) );
NAND3X1 NAND3X1_802 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_515_), .C(_516_), .Y(_517_) );
XNOR2X1 XNOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_2905_), .B(_328_), .Y(_518_) );
INVX1 INVX1_440 ( .gnd(gnd), .vdd(vdd), .A(_518_), .Y(_519_) );
NAND3X1 NAND3X1_803 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_517_), .C(_512_), .Y(_520_) );
AOI21X1 AOI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_516_), .C(_514_), .Y(_521_) );
AOI21X1 AOI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_511_), .C(_447_), .Y(_522_) );
OAI21X1 OAI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_522_), .C(_518_), .Y(_523_) );
NAND3X1 NAND3X1_804 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[37]), .B(_520_), .C(_523_), .Y(_524_) );
INVX1 INVX1_441 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[37]), .Y(_525_) );
NAND3X1 NAND3X1_805 ( .gnd(gnd), .vdd(vdd), .A(_518_), .B(_517_), .C(_512_), .Y(_526_) );
OAI21X1 OAI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_522_), .C(_519_), .Y(_527_) );
NAND3X1 NAND3X1_806 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(_526_), .C(_527_), .Y(_528_) );
NAND3X1 NAND3X1_807 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_524_), .C(_528_), .Y(_529_) );
NAND3X1 NAND3X1_808 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(_520_), .C(_523_), .Y(_530_) );
NAND3X1 NAND3X1_809 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[37]), .B(_526_), .C(_527_), .Y(_531_) );
NAND3X1 NAND3X1_810 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_530_), .C(_531_), .Y(_532_) );
NAND3X1 NAND3X1_811 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_532_), .C(_446_), .Y(_533_) );
INVX1 INVX1_442 ( .gnd(gnd), .vdd(vdd), .A(_9_), .Y(_534_) );
AOI21X1 AOI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_3689_), .C(_534_), .Y(_535_) );
NAND3X1 NAND3X1_812 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_530_), .C(_531_), .Y(_536_) );
NAND3X1 NAND3X1_813 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_524_), .C(_528_), .Y(_537_) );
NAND3X1 NAND3X1_814 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_536_), .C(_537_), .Y(_538_) );
XNOR2X1 XNOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_2970_), .B(_335_), .Y(_539_) );
INVX1 INVX1_443 ( .gnd(gnd), .vdd(vdd), .A(_539_), .Y(_540_) );
NAND3X1 NAND3X1_815 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_540_), .C(_533_), .Y(_541_) );
AOI21X1 AOI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_537_), .C(_535_), .Y(_542_) );
AOI21X1 AOI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_532_), .C(_446_), .Y(_543_) );
OAI21X1 OAI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_542_), .C(_539_), .Y(_544_) );
NAND3X1 NAND3X1_816 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[53]), .B(_541_), .C(_544_), .Y(_545_) );
INVX1 INVX1_444 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[53]), .Y(_546_) );
NAND3X1 NAND3X1_817 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_539_), .C(_533_), .Y(_547_) );
OAI21X1 OAI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_542_), .C(_540_), .Y(_548_) );
NAND3X1 NAND3X1_818 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(_547_), .C(_548_), .Y(_549_) );
NAND3X1 NAND3X1_819 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_545_), .C(_549_), .Y(_550_) );
NAND3X1 NAND3X1_820 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(_541_), .C(_544_), .Y(_551_) );
NAND3X1 NAND3X1_821 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[53]), .B(_547_), .C(_548_), .Y(_552_) );
NAND3X1 NAND3X1_822 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_551_), .C(_552_), .Y(_553_) );
NAND3X1 NAND3X1_823 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_550_), .C(_553_), .Y(_554_) );
AOI21X1 AOI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_36_), .C(_34_), .Y(_555_) );
AOI21X1 AOI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_3687_), .B(_37_), .C(_555_), .Y(_556_) );
NAND3X1 NAND3X1_824 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_551_), .C(_552_), .Y(_557_) );
NAND3X1 NAND3X1_825 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_545_), .C(_549_), .Y(_558_) );
NAND3X1 NAND3X1_826 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_557_), .C(_558_), .Y(_559_) );
XNOR2X1 XNOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_3058_), .B(_340_), .Y(_560_) );
INVX1 INVX1_445 ( .gnd(gnd), .vdd(vdd), .A(_560_), .Y(_561_) );
NAND3X1 NAND3X1_827 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_554_), .C(_559_), .Y(_562_) );
AOI21X1 AOI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_557_), .B(_558_), .C(_556_), .Y(_563_) );
AOI21X1 AOI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_553_), .C(_445_), .Y(_564_) );
OAI21X1 OAI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_564_), .C(_560_), .Y(_565_) );
NAND3X1 NAND3X1_828 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[69]), .B(_562_), .C(_565_), .Y(_566_) );
INVX1 INVX1_446 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[69]), .Y(_567_) );
NAND3X1 NAND3X1_829 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(_554_), .C(_559_), .Y(_568_) );
OAI21X1 OAI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_564_), .C(_561_), .Y(_569_) );
NAND3X1 NAND3X1_830 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_568_), .C(_569_), .Y(_570_) );
NAND3X1 NAND3X1_831 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_566_), .C(_570_), .Y(_571_) );
NAND3X1 NAND3X1_832 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_562_), .C(_565_), .Y(_572_) );
NAND3X1 NAND3X1_833 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[69]), .B(_568_), .C(_569_), .Y(_573_) );
NAND3X1 NAND3X1_834 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_572_), .C(_573_), .Y(_574_) );
NAND3X1 NAND3X1_835 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_571_), .C(_574_), .Y(_575_) );
AOI21X1 AOI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_60_), .C(_58_), .Y(_576_) );
AOI21X1 AOI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_3685_), .B(_61_), .C(_576_), .Y(_577_) );
NAND3X1 NAND3X1_836 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_572_), .C(_573_), .Y(_578_) );
NAND3X1 NAND3X1_837 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_566_), .C(_570_), .Y(_579_) );
NAND3X1 NAND3X1_838 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_578_), .C(_579_), .Y(_580_) );
NAND2X1 NAND2X1_430 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_344_), .Y(_581_) );
XNOR2X1 XNOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_3146_), .B(_581_), .Y(_582_) );
INVX1 INVX1_447 ( .gnd(gnd), .vdd(vdd), .A(_582_), .Y(_583_) );
NAND3X1 NAND3X1_839 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_580_), .C(_575_), .Y(_584_) );
AOI21X1 AOI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_578_), .B(_579_), .C(_577_), .Y(_585_) );
AOI21X1 AOI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_574_), .C(_443_), .Y(_586_) );
OAI21X1 OAI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_586_), .C(_582_), .Y(_587_) );
NAND3X1 NAND3X1_840 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[85]), .B(_584_), .C(_587_), .Y(_588_) );
INVX1 INVX1_448 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[85]), .Y(_589_) );
NAND3X1 NAND3X1_841 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_580_), .C(_575_), .Y(_590_) );
OAI21X1 OAI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_586_), .C(_583_), .Y(_591_) );
NAND3X1 NAND3X1_842 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_590_), .C(_591_), .Y(_592_) );
NAND3X1 NAND3X1_843 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_588_), .C(_592_), .Y(_593_) );
NAND3X1 NAND3X1_844 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_584_), .C(_587_), .Y(_594_) );
NAND3X1 NAND3X1_845 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[85]), .B(_590_), .C(_591_), .Y(_595_) );
NAND3X1 NAND3X1_846 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_594_), .C(_595_), .Y(_596_) );
NAND3X1 NAND3X1_847 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_596_), .C(_441_), .Y(_597_) );
AOI21X1 AOI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_84_), .C(_82_), .Y(_598_) );
AOI21X1 AOI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .B(_85_), .C(_598_), .Y(_599_) );
NAND3X1 NAND3X1_848 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_594_), .C(_595_), .Y(_600_) );
NAND3X1 NAND3X1_849 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_588_), .C(_592_), .Y(_601_) );
NAND3X1 NAND3X1_850 ( .gnd(gnd), .vdd(vdd), .A(_599_), .B(_600_), .C(_601_), .Y(_602_) );
XNOR2X1 XNOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_3190_), .B(_353_), .Y(_603_) );
NAND3X1 NAND3X1_851 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_602_), .C(_597_), .Y(_604_) );
AOI21X1 AOI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_601_), .C(_599_), .Y(_605_) );
AOI21X1 AOI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_596_), .C(_441_), .Y(_606_) );
INVX1 INVX1_449 ( .gnd(gnd), .vdd(vdd), .A(_603_), .Y(_607_) );
OAI21X1 OAI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_606_), .C(_607_), .Y(_608_) );
NAND3X1 NAND3X1_852 ( .gnd(gnd), .vdd(vdd), .A(W_133_), .B(_604_), .C(_608_), .Y(_609_) );
INVX1 INVX1_450 ( .gnd(gnd), .vdd(vdd), .A(W_133_), .Y(_610_) );
NAND3X1 NAND3X1_853 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_602_), .C(_597_), .Y(_611_) );
OAI21X1 OAI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_606_), .C(_603_), .Y(_612_) );
NAND3X1 NAND3X1_854 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_611_), .C(_612_), .Y(_613_) );
AOI21X1 AOI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_613_), .C(_104_), .Y(_614_) );
NAND3X1 NAND3X1_855 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_604_), .C(_608_), .Y(_615_) );
NAND3X1 NAND3X1_856 ( .gnd(gnd), .vdd(vdd), .A(W_133_), .B(_611_), .C(_612_), .Y(_616_) );
AOI21X1 AOI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_616_), .C(_108_), .Y(_617_) );
OAI21X1 OAI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_617_), .C(_439_), .Y(_618_) );
AOI21X1 AOI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_108_), .C(_106_), .Y(_619_) );
AOI21X1 AOI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_3680_), .B(_109_), .C(_619_), .Y(_620_) );
NAND3X1 NAND3X1_857 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_615_), .C(_616_), .Y(_621_) );
NAND3X1 NAND3X1_858 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_609_), .C(_613_), .Y(_622_) );
NAND3X1 NAND3X1_859 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_621_), .C(_622_), .Y(_623_) );
NAND3X1 NAND3X1_860 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_623_), .C(_618_), .Y(_624_) );
AOI21X1 AOI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_622_), .C(_620_), .Y(_625_) );
NAND3X1 NAND3X1_861 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_609_), .C(_613_), .Y(_626_) );
NAND3X1 NAND3X1_862 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_615_), .C(_616_), .Y(_627_) );
AOI21X1 AOI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_627_), .C(_439_), .Y(_628_) );
OAI21X1 OAI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_625_), .C(_360_), .Y(_629_) );
NAND2X1 NAND2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_629_), .Y(_630_) );
AOI21X1 AOI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_3198_), .B(_630_), .C(_437_), .Y(_631_) );
NAND3X1 NAND3X1_863 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_623_), .C(_618_), .Y(_632_) );
OAI21X1 OAI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_625_), .C(_361_), .Y(_633_) );
NAND3X1 NAND3X1_864 ( .gnd(gnd), .vdd(vdd), .A(_3198_), .B(_632_), .C(_633_), .Y(_634_) );
NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(W_149_), .B(_634_), .Y(_635_) );
OAI21X1 OAI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_631_), .C(_436_), .Y(_636_) );
NAND2X1 NAND2X1_432 ( .gnd(gnd), .vdd(vdd), .A(W_149_), .B(_634_), .Y(_637_) );
NAND3X1 NAND3X1_865 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_3198_), .C(_630_), .Y(_638_) );
NAND3X1 NAND3X1_866 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(_637_), .C(_638_), .Y(_639_) );
NAND3X1 NAND3X1_867 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_639_), .C(_636_), .Y(_640_) );
AOI21X1 AOI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_3677_), .B(_131_), .C(_134_), .Y(_641_) );
OAI21X1 OAI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_631_), .C(_123_), .Y(_642_) );
NAND3X1 NAND3X1_868 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_637_), .C(_638_), .Y(_643_) );
NAND3X1 NAND3X1_869 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_643_), .C(_642_), .Y(_644_) );
AOI21X1 AOI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_644_), .C(_369_), .Y(_645_) );
INVX1 INVX1_451 ( .gnd(gnd), .vdd(vdd), .A(_645_), .Y(_646_) );
NAND3X1 NAND3X1_870 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_640_), .C(_644_), .Y(_647_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_647_), .B(_3206_), .Y(_648_) );
AOI21X1 AOI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_646_), .B(_648_), .C(_434_), .Y(_649_) );
NAND2X1 NAND2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_3206_), .B(_647_), .Y(_650_) );
NOR3X1 NOR3X1_103 ( .gnd(gnd), .vdd(vdd), .A(W_165_), .B(_645_), .C(_650_), .Y(_651_) );
OAI21X1 OAI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_651_), .C(_433_), .Y(_652_) );
OAI21X1 OAI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_645_), .C(W_165_), .Y(_653_) );
NAND3X1 NAND3X1_871 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_646_), .C(_648_), .Y(_654_) );
NAND3X1 NAND3X1_872 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_653_), .C(_654_), .Y(_655_) );
NAND3X1 NAND3X1_873 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_655_), .C(_652_), .Y(_656_) );
AOI21X1 AOI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_3672_), .B(_155_), .C(_158_), .Y(_657_) );
OAI21X1 OAI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_651_), .C(_146_), .Y(_658_) );
NAND3X1 NAND3X1_874 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_653_), .C(_654_), .Y(_659_) );
NAND3X1 NAND3X1_875 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_659_), .C(_658_), .Y(_660_) );
NAND3X1 NAND3X1_876 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_656_), .C(_660_), .Y(_661_) );
AOI21X1 AOI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_658_), .C(_657_), .Y(_662_) );
AOI21X1 AOI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_652_), .C(_432_), .Y(_663_) );
OAI21X1 OAI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_663_), .C(_378_), .Y(_664_) );
NAND2X1 NAND2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_661_), .B(_664_), .Y(_665_) );
AOI21X1 AOI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_3214_), .B(_665_), .C(_431_), .Y(_666_) );
NAND3X1 NAND3X1_877 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_656_), .C(_660_), .Y(_667_) );
OAI21X1 OAI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_663_), .C(_380_), .Y(_668_) );
NAND3X1 NAND3X1_878 ( .gnd(gnd), .vdd(vdd), .A(_3214_), .B(_667_), .C(_668_), .Y(_669_) );
NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(W_181_), .B(_669_), .Y(_670_) );
OAI21X1 OAI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_666_), .C(_430_), .Y(_671_) );
NAND2X1 NAND2X1_435 ( .gnd(gnd), .vdd(vdd), .A(W_181_), .B(_669_), .Y(_672_) );
NAND3X1 NAND3X1_879 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_3214_), .C(_665_), .Y(_673_) );
NAND3X1 NAND3X1_880 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_672_), .C(_673_), .Y(_674_) );
NAND3X1 NAND3X1_881 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_429_), .C(_671_), .Y(_675_) );
AOI21X1 AOI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_3668_), .B(_179_), .C(_182_), .Y(_676_) );
OAI21X1 OAI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_666_), .C(_170_), .Y(_677_) );
NAND3X1 NAND3X1_882 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_672_), .C(_673_), .Y(_678_) );
NAND3X1 NAND3X1_883 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(_678_), .C(_677_), .Y(_679_) );
NAND3X1 NAND3X1_884 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_675_), .C(_679_), .Y(_680_) );
AOI21X1 AOI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_677_), .C(_676_), .Y(_681_) );
AOI21X1 AOI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_671_), .C(_429_), .Y(_682_) );
OAI21X1 OAI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_681_), .B(_682_), .C(_386_), .Y(_683_) );
NAND2X1 NAND2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(_683_), .Y(_684_) );
AOI21X1 AOI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .B(_684_), .C(_428_), .Y(_685_) );
NAND3X1 NAND3X1_885 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_675_), .C(_679_), .Y(_686_) );
OAI21X1 OAI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_681_), .B(_682_), .C(_388_), .Y(_687_) );
NAND3X1 NAND3X1_886 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .B(_686_), .C(_687_), .Y(_688_) );
NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(W_197_), .B(_688_), .Y(_689_) );
OAI21X1 OAI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_685_), .C(_427_), .Y(_690_) );
NAND2X1 NAND2X1_437 ( .gnd(gnd), .vdd(vdd), .A(W_197_), .B(_688_), .Y(_691_) );
NAND3X1 NAND3X1_887 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_3222_), .C(_684_), .Y(_692_) );
NAND3X1 NAND3X1_888 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_691_), .C(_692_), .Y(_693_) );
NAND3X1 NAND3X1_889 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_690_), .C(_426_), .Y(_694_) );
AOI21X1 AOI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_3663_), .B(_203_), .C(_206_), .Y(_695_) );
OAI21X1 OAI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_685_), .C(_194_), .Y(_696_) );
NAND3X1 NAND3X1_890 ( .gnd(gnd), .vdd(vdd), .A(_427_), .B(_691_), .C(_692_), .Y(_697_) );
NAND3X1 NAND3X1_891 ( .gnd(gnd), .vdd(vdd), .A(_697_), .B(_695_), .C(_696_), .Y(_698_) );
NAND3X1 NAND3X1_892 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_698_), .C(_694_), .Y(_699_) );
AOI21X1 AOI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_697_), .B(_696_), .C(_695_), .Y(_700_) );
AOI21X1 AOI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_690_), .C(_426_), .Y(_701_) );
OAI21X1 OAI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_701_), .C(_394_), .Y(_702_) );
NAND2X1 NAND2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_702_), .Y(_703_) );
AOI21X1 AOI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_3230_), .B(_703_), .C(_425_), .Y(_704_) );
NAND3X1 NAND3X1_893 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_698_), .C(_694_), .Y(_705_) );
OAI21X1 OAI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_701_), .C(_396_), .Y(_706_) );
NAND3X1 NAND3X1_894 ( .gnd(gnd), .vdd(vdd), .A(_3230_), .B(_705_), .C(_706_), .Y(_707_) );
NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(W_213_), .B(_707_), .Y(_708_) );
OAI21X1 OAI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_704_), .C(_424_), .Y(_709_) );
NAND2X1 NAND2X1_439 ( .gnd(gnd), .vdd(vdd), .A(W_213_), .B(_707_), .Y(_710_) );
NAND3X1 NAND3X1_895 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_3230_), .C(_703_), .Y(_711_) );
NAND3X1 NAND3X1_896 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_710_), .C(_711_), .Y(_712_) );
NAND3X1 NAND3X1_897 ( .gnd(gnd), .vdd(vdd), .A(_712_), .B(_423_), .C(_709_), .Y(_713_) );
AOI21X1 AOI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_3659_), .B(_229_), .C(_231_), .Y(_714_) );
OAI21X1 OAI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_704_), .C(_220_), .Y(_715_) );
NAND3X1 NAND3X1_898 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_710_), .C(_711_), .Y(_716_) );
NAND3X1 NAND3X1_899 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_716_), .C(_715_), .Y(_717_) );
NAND3X1 NAND3X1_900 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_713_), .C(_717_), .Y(_718_) );
AOI21X1 AOI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_715_), .C(_714_), .Y(_719_) );
AOI21X1 AOI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_712_), .B(_709_), .C(_423_), .Y(_720_) );
OAI21X1 OAI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_720_), .C(_402_), .Y(_721_) );
NAND2X1 NAND2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_721_), .Y(_722_) );
AOI21X1 AOI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_3238_), .B(_722_), .C(_422_), .Y(_723_) );
NAND3X1 NAND3X1_901 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_713_), .C(_717_), .Y(_724_) );
OAI21X1 OAI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_720_), .C(_404_), .Y(_725_) );
NAND3X1 NAND3X1_902 ( .gnd(gnd), .vdd(vdd), .A(_3238_), .B(_724_), .C(_725_), .Y(_726_) );
NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(W_229_), .B(_726_), .Y(_727_) );
OAI21X1 OAI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_723_), .C(_421_), .Y(_728_) );
NAND2X1 NAND2X1_441 ( .gnd(gnd), .vdd(vdd), .A(W_229_), .B(_726_), .Y(_729_) );
NAND3X1 NAND3X1_903 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(_3238_), .C(_722_), .Y(_730_) );
NAND3X1 NAND3X1_904 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_729_), .C(_730_), .Y(_731_) );
NAND3X1 NAND3X1_905 ( .gnd(gnd), .vdd(vdd), .A(_420_), .B(_731_), .C(_728_), .Y(_732_) );
AOI21X1 AOI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_3653_), .C(_256_), .Y(_733_) );
OAI21X1 OAI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_723_), .C(_245_), .Y(_734_) );
NAND3X1 NAND3X1_906 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_729_), .C(_730_), .Y(_735_) );
NAND3X1 NAND3X1_907 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_733_), .C(_734_), .Y(_736_) );
AOI21X1 AOI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_736_), .C(_410_), .Y(_737_) );
NAND3X1 NAND3X1_908 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_732_), .C(_736_), .Y(_738_) );
NAND2X1 NAND2X1_442 ( .gnd(gnd), .vdd(vdd), .A(_3247_), .B(_738_), .Y(_739_) );
OAI21X1 OAI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(_739_), .B(_737_), .C(W_245_), .Y(_740_) );
INVX1 INVX1_452 ( .gnd(gnd), .vdd(vdd), .A(W_245_), .Y(_741_) );
INVX1 INVX1_453 ( .gnd(gnd), .vdd(vdd), .A(_737_), .Y(_742_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_738_), .B(_3247_), .Y(_743_) );
NAND3X1 NAND3X1_909 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_742_), .C(_743_), .Y(_744_) );
AOI21X1 AOI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_740_), .B(_744_), .C(_268_), .Y(_745_) );
INVX1 INVX1_454 ( .gnd(gnd), .vdd(vdd), .A(_268_), .Y(_746_) );
AOI21X1 AOI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_742_), .B(_743_), .C(_741_), .Y(_747_) );
NOR3X1 NOR3X1_104 ( .gnd(gnd), .vdd(vdd), .A(W_245_), .B(_737_), .C(_739_), .Y(_748_) );
NOR3X1 NOR3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_748_), .C(_747_), .Y(_749_) );
OAI21X1 OAI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_745_), .C(_419_), .Y(_750_) );
AOI21X1 AOI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_3651_), .C(_281_), .Y(_751_) );
OAI21X1 OAI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_748_), .C(_746_), .Y(_752_) );
NAND3X1 NAND3X1_910 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_740_), .C(_744_), .Y(_753_) );
NAND3X1 NAND3X1_911 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_752_), .C(_751_), .Y(_754_) );
NAND3X1 NAND3X1_912 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_754_), .C(_750_), .Y(_755_) );
NAND3X1 NAND3X1_913 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_419_), .C(_752_), .Y(_756_) );
OAI21X1 OAI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_745_), .C(_751_), .Y(_757_) );
NAND3X1 NAND3X1_914 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_756_), .C(_757_), .Y(_758_) );
AOI21X1 AOI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_758_), .C(_292_), .Y(_759_) );
NAND2X1 NAND2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_758_), .Y(_760_) );
NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_760_), .Y(_761_) );
NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_761_), .Y(H_5_) );
OAI21X1 OAI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_751_), .C(_752_), .Y(_762_) );
AOI21X1 AOI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_730_), .C(_245_), .Y(_763_) );
AOI21X1 AOI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_420_), .B(_731_), .C(_763_), .Y(_764_) );
INVX2 INVX2_138 ( .gnd(gnd), .vdd(vdd), .A(W_230_), .Y(_765_) );
NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_3446_), .B(_3443_), .Y(_766_) );
INVX2 INVX2_139 ( .gnd(gnd), .vdd(vdd), .A(_766_), .Y(_767_) );
AOI21X1 AOI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_710_), .B(_711_), .C(_220_), .Y(_768_) );
AOI21X1 AOI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_712_), .B(_423_), .C(_768_), .Y(_769_) );
INVX2 INVX2_140 ( .gnd(gnd), .vdd(vdd), .A(W_214_), .Y(_770_) );
AOI21X1 AOI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_691_), .B(_692_), .C(_194_), .Y(_771_) );
AOI21X1 AOI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_426_), .C(_771_), .Y(_772_) );
INVX2 INVX2_141 ( .gnd(gnd), .vdd(vdd), .A(W_198_), .Y(_773_) );
NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_3419_), .B(_3416_), .Y(_774_) );
INVX2 INVX2_142 ( .gnd(gnd), .vdd(vdd), .A(_774_), .Y(_775_) );
AOI21X1 AOI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_673_), .C(_170_), .Y(_776_) );
AOI21X1 AOI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_429_), .C(_776_), .Y(_777_) );
INVX2 INVX2_143 ( .gnd(gnd), .vdd(vdd), .A(W_182_), .Y(_778_) );
NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_3407_), .B(_3405_), .Y(_779_) );
INVX2 INVX2_144 ( .gnd(gnd), .vdd(vdd), .A(_779_), .Y(_780_) );
INVX1 INVX1_455 ( .gnd(gnd), .vdd(vdd), .A(_652_), .Y(_781_) );
AOI21X1 AOI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_432_), .C(_781_), .Y(_782_) );
INVX2 INVX2_145 ( .gnd(gnd), .vdd(vdd), .A(W_166_), .Y(_783_) );
NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .B(_3396_), .Y(_784_) );
INVX1 INVX1_456 ( .gnd(gnd), .vdd(vdd), .A(_784_), .Y(_785_) );
INVX1 INVX1_457 ( .gnd(gnd), .vdd(vdd), .A(_636_), .Y(_786_) );
AOI21X1 AOI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_639_), .C(_786_), .Y(_787_) );
INVX2 INVX2_146 ( .gnd(gnd), .vdd(vdd), .A(W_150_), .Y(_788_) );
NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_3381_), .B(_3383_), .Y(_789_) );
INVX1 INVX1_458 ( .gnd(gnd), .vdd(vdd), .A(_789_), .Y(_790_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_626_), .Y(_791_) );
INVX1 INVX1_459 ( .gnd(gnd), .vdd(vdd), .A(W_134_), .Y(_792_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_597_), .B(_593_), .Y(_793_) );
INVX1 INVX1_460 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[86]), .Y(_794_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_571_), .Y(_795_) );
INVX1 INVX1_461 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[70]), .Y(_796_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_550_), .Y(_797_) );
INVX1 INVX1_462 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[54]), .Y(_798_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_529_), .Y(_799_) );
INVX1 INVX1_463 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[38]), .Y(_800_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_508_), .Y(_801_) );
INVX1 INVX1_464 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[22]), .Y(_802_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_493_), .Y(_803_) );
INVX1 INVX1_465 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[6]), .Y(_804_) );
OAI21X1 OAI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_474_), .C(_472_), .Y(_805_) );
INVX2 INVX2_147 ( .gnd(gnd), .vdd(vdd), .A(_805_), .Y(_806_) );
INVX1 INVX1_466 ( .gnd(gnd), .vdd(vdd), .A(_466_), .Y(_807_) );
INVX1 INVX1_467 ( .gnd(gnd), .vdd(vdd), .A(W_22_), .Y(_808_) );
NAND2X1 NAND2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_3288_), .B(_3292_), .Y(_809_) );
XNOR2X1 XNOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(W_6_), .Y(_810_) );
XNOR2X1 XNOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_810_), .B(_809_), .Y(_811_) );
NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_808_), .B(_811_), .Y(_812_) );
XOR2X1 XOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_810_), .B(_809_), .Y(_813_) );
NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(W_22_), .B(_813_), .Y(_814_) );
NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_814_), .Y(_815_) );
NAND2X1 NAND2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_807_), .B(_815_), .Y(_816_) );
OAI21X1 OAI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_814_), .B(_812_), .C(_466_), .Y(_817_) );
NAND2X1 NAND2X1_446 ( .gnd(gnd), .vdd(vdd), .A(_817_), .B(_816_), .Y(_818_) );
NAND2X1 NAND2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_806_), .B(_818_), .Y(_819_) );
XNOR2X1 XNOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_815_), .B(_466_), .Y(_820_) );
NAND2X1 NAND2X1_448 ( .gnd(gnd), .vdd(vdd), .A(_805_), .B(_820_), .Y(_821_) );
INVX2 INVX2_148 ( .gnd(gnd), .vdd(vdd), .A(W_10_), .Y(_822_) );
NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_3299_), .B(_3303_), .Y(_823_) );
XNOR2X1 XNOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_823_), .B(_822_), .Y(_824_) );
NAND3X1 NAND3X1_915 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(_819_), .C(_821_), .Y(_825_) );
NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_805_), .B(_820_), .Y(_826_) );
NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_806_), .B(_818_), .Y(_827_) );
INVX1 INVX1_468 ( .gnd(gnd), .vdd(vdd), .A(_824_), .Y(_828_) );
OAI21X1 OAI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_826_), .B(_827_), .C(_828_), .Y(_829_) );
NAND3X1 NAND3X1_916 ( .gnd(gnd), .vdd(vdd), .A(_804_), .B(_825_), .C(_829_), .Y(_830_) );
NAND3X1 NAND3X1_917 ( .gnd(gnd), .vdd(vdd), .A(_828_), .B(_819_), .C(_821_), .Y(_831_) );
OAI21X1 OAI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(_826_), .B(_827_), .C(_824_), .Y(_832_) );
NAND3X1 NAND3X1_918 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[6]), .B(_831_), .C(_832_), .Y(_833_) );
AOI21X1 AOI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_830_), .B(_833_), .C(_488_), .Y(_834_) );
INVX1 INVX1_469 ( .gnd(gnd), .vdd(vdd), .A(_488_), .Y(_835_) );
NAND3X1 NAND3X1_919 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[6]), .B(_825_), .C(_829_), .Y(_836_) );
NAND3X1 NAND3X1_920 ( .gnd(gnd), .vdd(vdd), .A(_804_), .B(_831_), .C(_832_), .Y(_837_) );
AOI21X1 AOI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_836_), .B(_837_), .C(_835_), .Y(_838_) );
OAI21X1 OAI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_834_), .B(_838_), .C(_803_), .Y(_839_) );
NAND2X1 NAND2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_499_), .Y(_840_) );
NAND3X1 NAND3X1_921 ( .gnd(gnd), .vdd(vdd), .A(_835_), .B(_836_), .C(_837_), .Y(_841_) );
NAND3X1 NAND3X1_922 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_830_), .C(_833_), .Y(_842_) );
NAND3X1 NAND3X1_923 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_841_), .C(_842_), .Y(_843_) );
NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_3310_), .B(_3313_), .Y(_844_) );
OAI21X1 OAI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(W_24_), .B(W_8_), .C(_316_), .Y(_845_) );
INVX1 INVX1_470 ( .gnd(gnd), .vdd(vdd), .A(W_26_), .Y(_846_) );
NAND2X1 NAND2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_822_), .Y(_847_) );
NAND2X1 NAND2X1_451 ( .gnd(gnd), .vdd(vdd), .A(W_26_), .B(W_10_), .Y(_848_) );
NAND2X1 NAND2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_847_), .Y(_849_) );
OAI21X1 OAI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_314_), .C(_849_), .Y(_850_) );
NAND3X1 NAND3X1_924 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_848_), .C(_315_), .Y(_851_) );
NAND2X1 NAND2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_851_), .B(_850_), .Y(_852_) );
NAND2X1 NAND2X1_454 ( .gnd(gnd), .vdd(vdd), .A(_845_), .B(_852_), .Y(_853_) );
NAND3X1 NAND3X1_925 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_851_), .C(_317_), .Y(_854_) );
NAND2X1 NAND2X1_455 ( .gnd(gnd), .vdd(vdd), .A(_854_), .B(_853_), .Y(_855_) );
XNOR2X1 XNOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_855_), .Y(_856_) );
NAND3X1 NAND3X1_926 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_856_), .C(_839_), .Y(_857_) );
AOI21X1 AOI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_841_), .B(_842_), .C(_840_), .Y(_858_) );
NOR3X1 NOR3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_834_), .B(_838_), .C(_803_), .Y(_859_) );
INVX1 INVX1_471 ( .gnd(gnd), .vdd(vdd), .A(_856_), .Y(_860_) );
OAI21X1 OAI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(_858_), .C(_860_), .Y(_861_) );
NAND3X1 NAND3X1_927 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_857_), .C(_861_), .Y(_862_) );
NAND3X1 NAND3X1_928 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_860_), .C(_839_), .Y(_863_) );
OAI21X1 OAI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(_858_), .C(_856_), .Y(_864_) );
NAND3X1 NAND3X1_929 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[22]), .B(_863_), .C(_864_), .Y(_865_) );
AOI21X1 AOI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_865_), .C(_503_), .Y(_866_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(_3860_) );
NAND2X1 NAND2X1_456 ( .gnd(gnd), .vdd(vdd), .A(W_1_), .B(W_0_), .Y(_3861_) );
NAND2X1 NAND2X1_457 ( .gnd(gnd), .vdd(vdd), .A(W_3_), .B(W_2_), .Y(_3862_) );
NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_3861_), .B(_3862_), .Y(_3863_) );
NAND2X1 NAND2X1_458 ( .gnd(gnd), .vdd(vdd), .A(W_6_), .B(W_5_), .Y(_3864_) );
NAND2X1 NAND2X1_459 ( .gnd(gnd), .vdd(vdd), .A(W_7_), .B(W_4_), .Y(_3865_) );
NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_3864_), .B(_3865_), .Y(_3866_) );
NAND2X1 NAND2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_3863_), .B(_3866_), .Y(_3867_) );
NAND2X1 NAND2X1_461 ( .gnd(gnd), .vdd(vdd), .A(W_10_), .B(W_9_), .Y(_3868_) );
NAND2X1 NAND2X1_462 ( .gnd(gnd), .vdd(vdd), .A(W_11_), .B(W_8_), .Y(_3869_) );
NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_3868_), .B(_3869_), .Y(_3870_) );
NAND2X1 NAND2X1_463 ( .gnd(gnd), .vdd(vdd), .A(W_14_), .B(W_13_), .Y(_3871_) );
NAND2X1 NAND2X1_464 ( .gnd(gnd), .vdd(vdd), .A(W_15_), .B(W_12_), .Y(_3872_) );
NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_3872_), .Y(_3873_) );
NAND2X1 NAND2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_3870_), .B(_3873_), .Y(_3874_) );
NAND2X1 NAND2X1_466 ( .gnd(gnd), .vdd(vdd), .A(W_18_), .B(W_17_), .Y(_3875_) );
NAND2X1 NAND2X1_467 ( .gnd(gnd), .vdd(vdd), .A(W_19_), .B(W_16_), .Y(_3876_) );
NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_3875_), .B(_3876_), .Y(_3877_) );
INVX1 INVX1_472 ( .gnd(gnd), .vdd(vdd), .A(_3877_), .Y(_3878_) );
NOR3X1 NOR3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_3867_), .B(_3878_), .C(_3874_), .Y(_3879_) );
INVX1 INVX1_473 ( .gnd(gnd), .vdd(vdd), .A(W_26_), .Y(_3880_) );
INVX2 INVX2_149 ( .gnd(gnd), .vdd(vdd), .A(W_25_), .Y(_3881_) );
NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_3880_), .B(_3881_), .Y(_3882_) );
INVX2 INVX2_150 ( .gnd(gnd), .vdd(vdd), .A(_3882_), .Y(_3883_) );
NAND2X1 NAND2X1_468 ( .gnd(gnd), .vdd(vdd), .A(W_27_), .B(W_24_), .Y(_3884_) );
NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_3884_), .B(_3883_), .Y(_3885_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(W_29_), .Y(_3886_) );
INVX1 INVX1_474 ( .gnd(gnd), .vdd(vdd), .A(W_28_), .Y(_3887_) );
NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_3886_), .B(_3887_), .Y(_3888_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(W_23_), .B(W_20_), .Y(_3889_) );
NAND2X1 NAND2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_3889_), .B(_3888_), .Y(_3890_) );
INVX1 INVX1_475 ( .gnd(gnd), .vdd(vdd), .A(W_31_), .Y(_3891_) );
INVX2 INVX2_151 ( .gnd(gnd), .vdd(vdd), .A(W_30_), .Y(_3892_) );
NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_3891_), .B(_3892_), .Y(_3893_) );
NAND2X1 NAND2X1_470 ( .gnd(gnd), .vdd(vdd), .A(W_22_), .B(W_21_), .Y(_3773_) );
INVX1 INVX1_476 ( .gnd(gnd), .vdd(vdd), .A(_3773_), .Y(_3774_) );
NAND2X1 NAND2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_3774_), .B(_3893_), .Y(_3775_) );
NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_3890_), .B(_3775_), .Y(_3776_) );
NAND3X1 NAND3X1_930 ( .gnd(gnd), .vdd(vdd), .A(_3885_), .B(_3776_), .C(_3879_), .Y(_3777_) );
AOI21X1 AOI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(W_0_), .B(_3777__bF_buf4), .C(_3860__bF_buf4), .Y(_3772__0_) );
XNOR2X1 XNOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(W_1_), .B(W_0_), .Y(_3778_) );
AOI21X1 AOI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_3778_), .B(_3777__bF_buf1), .C(_3860__bF_buf1), .Y(_3772__1_) );
XOR2X1 XOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_3861_), .B(W_2_), .Y(_3779_) );
AOI21X1 AOI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_3779_), .B(_3777__bF_buf1), .C(_3860__bF_buf1), .Y(_3772__2_) );
INVX1 INVX1_477 ( .gnd(gnd), .vdd(vdd), .A(_3863_), .Y(_3780_) );
NAND3X1 NAND3X1_931 ( .gnd(gnd), .vdd(vdd), .A(W_2_), .B(W_1_), .C(W_0_), .Y(_3781_) );
INVX1 INVX1_478 ( .gnd(gnd), .vdd(vdd), .A(_3781_), .Y(_3782_) );
OAI21X1 OAI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_3782_), .B(W_3_), .C(_3780_), .Y(_3783_) );
AOI21X1 AOI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_3783_), .B(_3777__bF_buf1), .C(_3860__bF_buf1), .Y(_3772__3_) );
XNOR2X1 XNOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_3863_), .B(W_4_), .Y(_3784_) );
AOI21X1 AOI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_3784_), .B(_3777__bF_buf0), .C(_3860__bF_buf3), .Y(_3772__4_) );
INVX1 INVX1_479 ( .gnd(gnd), .vdd(vdd), .A(W_5_), .Y(_3785_) );
NAND2X1 NAND2X1_472 ( .gnd(gnd), .vdd(vdd), .A(W_4_), .B(_3863_), .Y(_3786_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_3786_), .B(_3785_), .Y(_3787_) );
NAND2X1 NAND2X1_473 ( .gnd(gnd), .vdd(vdd), .A(_3785_), .B(_3786_), .Y(_3788_) );
NAND2X1 NAND2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_3788_), .B(_3787_), .Y(_3789_) );
AOI21X1 AOI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_3789_), .B(_3777__bF_buf0), .C(_3860__bF_buf3), .Y(_3772__5_) );
XOR2X1 XOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_3787_), .B(W_6_), .Y(_3790_) );
AOI21X1 AOI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf0), .B(_3790_), .C(_3860__bF_buf3), .Y(_3772__6_) );
NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_3864_), .B(_3786_), .Y(_3791_) );
OAI21X1 OAI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_3791_), .B(W_7_), .C(_3867_), .Y(_3792_) );
AOI21X1 AOI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_3792_), .B(_3777__bF_buf1), .C(_3860__bF_buf1), .Y(_3772__7_) );
INVX1 INVX1_480 ( .gnd(gnd), .vdd(vdd), .A(W_8_), .Y(_3793_) );
NAND2X1 NAND2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_3793_), .B(_3867_), .Y(_3794_) );
INVX1 INVX1_481 ( .gnd(gnd), .vdd(vdd), .A(_3867_), .Y(_3795_) );
NAND2X1 NAND2X1_476 ( .gnd(gnd), .vdd(vdd), .A(W_8_), .B(_3795_), .Y(_3796_) );
NAND2X1 NAND2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_3794_), .B(_3796_), .Y(_3797_) );
AOI21X1 AOI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_3797_), .B(_3777__bF_buf0), .C(_3860__bF_buf3), .Y(_3772__8_) );
INVX2 INVX2_152 ( .gnd(gnd), .vdd(vdd), .A(W_9_), .Y(_3798_) );
XNOR2X1 XNOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_3796_), .B(_3798_), .Y(_3799_) );
AOI21X1 AOI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf0), .B(_3799_), .C(_3860__bF_buf3), .Y(_3772__9_) );
INVX1 INVX1_482 ( .gnd(gnd), .vdd(vdd), .A(W_10_), .Y(_3800_) );
OAI21X1 OAI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_3796_), .B(_3798_), .C(_3800_), .Y(_3801_) );
OAI21X1 OAI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_3868_), .B(_3796_), .C(_3801_), .Y(_3802_) );
AOI21X1 AOI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf0), .B(_3802_), .C(_3860__bF_buf3), .Y(_3772__10_) );
NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_3868_), .B(_3796_), .Y(_3803_) );
NAND2X1 NAND2X1_478 ( .gnd(gnd), .vdd(vdd), .A(_3870_), .B(_3795_), .Y(_3804_) );
OAI21X1 OAI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_3803_), .B(W_11_), .C(_3804_), .Y(_3805_) );
AOI21X1 AOI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf3), .B(_3805_), .C(_3860__bF_buf0), .Y(_3772__11_) );
INVX1 INVX1_483 ( .gnd(gnd), .vdd(vdd), .A(W_12_), .Y(_3806_) );
NAND2X1 NAND2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_3806_), .B(_3804_), .Y(_3807_) );
OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_3804_), .B(_3806_), .Y(_3808_) );
NAND2X1 NAND2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_3807_), .B(_3808_), .Y(_3809_) );
AOI21X1 AOI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf3), .B(_3809_), .C(_3860__bF_buf0), .Y(_3772__12_) );
INVX2 INVX2_153 ( .gnd(gnd), .vdd(vdd), .A(W_13_), .Y(_3810_) );
XNOR2X1 XNOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3808_), .B(_3810_), .Y(_3811_) );
AOI21X1 AOI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf3), .B(_3811_), .C(_3860__bF_buf0), .Y(_3772__13_) );
INVX1 INVX1_484 ( .gnd(gnd), .vdd(vdd), .A(W_14_), .Y(_3812_) );
OAI21X1 OAI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_3808_), .B(_3810_), .C(_3812_), .Y(_3813_) );
OAI21X1 OAI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_3808_), .C(_3813_), .Y(_3814_) );
AOI21X1 AOI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf3), .B(_3814_), .C(_3860__bF_buf0), .Y(_3772__14_) );
NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_3867_), .B(_3874_), .Y(_3815_) );
INVX1 INVX1_485 ( .gnd(gnd), .vdd(vdd), .A(_3815_), .Y(_3816_) );
NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_3808_), .Y(_3817_) );
OAI21X1 OAI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_3817_), .B(W_15_), .C(_3816_), .Y(_3818_) );
AOI21X1 AOI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf3), .B(_3818_), .C(_3860__bF_buf0), .Y(_3772__15_) );
XNOR2X1 XNOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_3815_), .B(W_16_), .Y(_3819_) );
AOI21X1 AOI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf3), .B(_3819_), .C(_3860__bF_buf0), .Y(_3772__16_) );
INVX2 INVX2_154 ( .gnd(gnd), .vdd(vdd), .A(W_17_), .Y(_3820_) );
NAND2X1 NAND2X1_481 ( .gnd(gnd), .vdd(vdd), .A(W_16_), .B(_3815_), .Y(_3821_) );
XNOR2X1 XNOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_3821_), .B(_3820_), .Y(_3822_) );
AOI21X1 AOI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf4), .B(_3822_), .C(_3860__bF_buf4), .Y(_3772__17_) );
INVX1 INVX1_486 ( .gnd(gnd), .vdd(vdd), .A(W_18_), .Y(_3823_) );
OAI21X1 OAI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_3821_), .B(_3820_), .C(_3823_), .Y(_3824_) );
OAI21X1 OAI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_3875_), .B(_3821_), .C(_3824_), .Y(_3825_) );
AOI21X1 AOI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf4), .B(_3825_), .C(_3860__bF_buf4), .Y(_3772__18_) );
INVX1 INVX1_487 ( .gnd(gnd), .vdd(vdd), .A(_3879_), .Y(_3826_) );
NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_3875_), .B(_3821_), .Y(_3827_) );
OAI21X1 OAI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_3827_), .B(W_19_), .C(_3826_), .Y(_3828_) );
AOI21X1 AOI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf4), .B(_3828_), .C(_3860__bF_buf4), .Y(_3772__19_) );
NAND3X1 NAND3X1_932 ( .gnd(gnd), .vdd(vdd), .A(W_20_), .B(_3877_), .C(_3815_), .Y(_3829_) );
AOI21X1 AOI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_3885_), .B(_3776_), .C(_3829_), .Y(_3830_) );
OAI21X1 OAI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_3879_), .B(W_20_), .C(inicio), .Y(_3831_) );
NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_3831_), .B(_3830_), .Y(_3772__20_) );
INVX2 INVX2_155 ( .gnd(gnd), .vdd(vdd), .A(W_21_), .Y(_3832_) );
XNOR2X1 XNOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_3829_), .B(_3832_), .Y(_3833_) );
AOI21X1 AOI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf4), .B(_3833_), .C(_3860__bF_buf4), .Y(_3772__21_) );
NOR2X1 NOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_3832_), .B(_3829_), .Y(_3834_) );
NAND3X1 NAND3X1_933 ( .gnd(gnd), .vdd(vdd), .A(W_20_), .B(_3774_), .C(_3879_), .Y(_3835_) );
OAI21X1 OAI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_3834_), .B(W_22_), .C(_3835_), .Y(_3836_) );
AOI21X1 AOI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf2), .B(_3836_), .C(_3860__bF_buf2), .Y(_3772__22_) );
INVX2 INVX2_156 ( .gnd(gnd), .vdd(vdd), .A(W_23_), .Y(_3837_) );
OAI21X1 OAI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_3829_), .B(_3773_), .C(_3837_), .Y(_3838_) );
NOR3X1 NOR3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_3837_), .B(_3773_), .C(_3829_), .Y(_3839_) );
INVX1 INVX1_488 ( .gnd(gnd), .vdd(vdd), .A(_3839_), .Y(_3840_) );
NAND2X1 NAND2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_3838_), .B(_3840_), .Y(_3841_) );
AOI21X1 AOI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf2), .B(_3841_), .C(_3860__bF_buf2), .Y(_3772__23_) );
XNOR2X1 XNOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_3839_), .B(W_24_), .Y(_3842_) );
AOI21X1 AOI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf2), .B(_3842_), .C(_3860__bF_buf2), .Y(_3772__24_) );
NAND2X1 NAND2X1_483 ( .gnd(gnd), .vdd(vdd), .A(W_24_), .B(_3839_), .Y(_3843_) );
XNOR2X1 XNOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_3843_), .B(_3881_), .Y(_3844_) );
AOI21X1 AOI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf4), .B(_3844_), .C(_3860__bF_buf4), .Y(_3772__25_) );
OAI21X1 OAI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_3843_), .B(_3881_), .C(_3880_), .Y(_3845_) );
OAI21X1 OAI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_3883_), .B(_3843_), .C(_3845_), .Y(_3846_) );
AOI21X1 AOI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf2), .B(_3846_), .C(_3860__bF_buf4), .Y(_3772__26_) );
NOR2X1 NOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_3883_), .B(_3843_), .Y(_3847_) );
INVX1 INVX1_489 ( .gnd(gnd), .vdd(vdd), .A(_3885_), .Y(_3848_) );
NOR3X1 NOR3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_3837_), .B(_3848_), .C(_3835_), .Y(_3849_) );
INVX1 INVX1_490 ( .gnd(gnd), .vdd(vdd), .A(_3849_), .Y(_3850_) );
OAI21X1 OAI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_3847_), .B(W_27_), .C(_3850_), .Y(_3851_) );
AOI21X1 AOI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf2), .B(_3851_), .C(_3860__bF_buf2), .Y(_3772__27_) );
OAI21X1 OAI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_3840_), .B(_3848_), .C(_3887_), .Y(_3852_) );
NAND3X1 NAND3X1_934 ( .gnd(gnd), .vdd(vdd), .A(W_28_), .B(_3885_), .C(_3839_), .Y(_3853_) );
NAND2X1 NAND2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(_3852_), .Y(_3854_) );
AOI21X1 AOI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf2), .B(_3854_), .C(_3860__bF_buf2), .Y(_3772__28_) );
XNOR2X1 XNOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(_3886_), .Y(_3855_) );
AOI21X1 AOI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf1), .B(_3855_), .C(_3860__bF_buf2), .Y(_3772__29_) );
OAI21X1 OAI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(_3886_), .C(_3892_), .Y(_3856_) );
NOR2X1 NOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_3892_), .B(_3886_), .Y(_3857_) );
NAND3X1 NAND3X1_935 ( .gnd(gnd), .vdd(vdd), .A(W_28_), .B(_3857_), .C(_3849_), .Y(_3858_) );
NAND2X1 NAND2X1_485 ( .gnd(gnd), .vdd(vdd), .A(_3858_), .B(_3856_), .Y(_3859_) );
AOI21X1 AOI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_3777__bF_buf1), .B(_3859_), .C(_3860__bF_buf1), .Y(_3772__30_) );
AOI21X1 AOI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_3891_), .B(_3858_), .C(_3860__bF_buf1), .Y(_3772__31_) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3772__0_), .Q(W_0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3772__1_), .Q(W_1_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3772__2_), .Q(W_2_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3772__3_), .Q(W_3_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3772__4_), .Q(W_4_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3772__5_), .Q(W_5_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3772__6_), .Q(W_6_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3772__7_), .Q(W_7_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3772__8_), .Q(W_8_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3772__9_), .Q(W_9_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3772__10_), .Q(W_10_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3772__11_), .Q(W_11_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3772__12_), .Q(W_12_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3772__13_), .Q(W_13_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3772__14_), .Q(W_14_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3772__15_), .Q(W_15_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3772__16_), .Q(W_16_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3772__17_), .Q(W_17_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3772__18_), .Q(W_18_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3772__19_), .Q(W_19_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3772__20_), .Q(W_20_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3772__21_), .Q(W_21_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3772__22_), .Q(W_22_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3772__23_), .Q(W_23_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3772__24_), .Q(W_24_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3772__25_), .Q(W_25_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3772__26_), .Q(W_26_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3772__27_), .Q(W_27_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3772__28_), .Q(W_28_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3772__29_), .Q(W_29_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3772__30_), .Q(W_30_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3772__31_), .Q(W_31_) );
INVX1 INVX1_491 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_3931_) );
INVX1 INVX1_492 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .Y(_3932_) );
INVX1 INVX1_493 ( .gnd(gnd), .vdd(vdd), .A(target[0]), .Y(_3933_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3932_), .B(gnd), .C(_3933_), .D(vdd), .Y(_3934_) );
OAI21X1 OAI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .B(_3931_), .C(_3934_), .Y(_3935_) );
XOR2X1 XOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(vdd), .Y(_3936_) );
INVX2 INVX2_157 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .Y(_3937_) );
INVX1 INVX1_494 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_3938_) );
NAND2X1 NAND2X1_486 ( .gnd(gnd), .vdd(vdd), .A(_3937_), .B(_3938_), .Y(_3939_) );
NAND2X1 NAND2X1_487 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(gnd), .Y(_3940_) );
AOI21X1 AOI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_3939_), .B(_3940_), .C(_3936_), .Y(_3941_) );
INVX1 INVX1_495 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .Y(_3942_) );
NAND2X1 NAND2X1_488 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_3942_), .Y(_3943_) );
NAND2X1 NAND2X1_489 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_3937_), .Y(_3944_) );
OAI21X1 OAI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_3936_), .B(_3944_), .C(_3943_), .Y(_3945_) );
AOI21X1 AOI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_3941_), .C(_3945_), .Y(_3946_) );
INVX1 INVX1_496 ( .gnd(gnd), .vdd(vdd), .A(H_15_), .Y(_3947_) );
INVX1 INVX1_497 ( .gnd(gnd), .vdd(vdd), .A(H_14_), .Y(_3948_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_3947_), .B(target[7]), .C(target[6]), .D(_3948_), .Y(_3949_) );
INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .Y(_3950_) );
INVX2 INVX2_158 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .Y(_3951_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_3950_), .B(H_15_), .C(_3951_), .D(H_14_), .Y(_3952_) );
NOR2X1 NOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_3949_), .B(_3952_), .Y(_3953_) );
INVX2 INVX2_159 ( .gnd(gnd), .vdd(vdd), .A(H_13_), .Y(_3954_) );
INVX1 INVX1_498 ( .gnd(gnd), .vdd(vdd), .A(H_12_), .Y(_3955_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_3954_), .B(target[5]), .C(target[4]), .D(_3955_), .Y(_3956_) );
INVX2 INVX2_160 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .Y(_3957_) );
INVX1 INVX1_499 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .Y(_3958_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_3957_), .B(H_13_), .C(_3958_), .D(H_12_), .Y(_3959_) );
NOR2X1 NOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_3956_), .B(_3959_), .Y(_3960_) );
NAND2X1 NAND2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_3953_), .B(_3960_), .Y(_3961_) );
NAND2X1 NAND2X1_491 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .B(_3954_), .Y(_3962_) );
NAND3X1 NAND3X1_936 ( .gnd(gnd), .vdd(vdd), .A(_3956_), .B(_3962_), .C(_3953_), .Y(_3963_) );
OAI21X1 OAI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_3946_), .B(_3961_), .C(_3963_), .Y(_3964_) );
INVX1 INVX1_500 ( .gnd(gnd), .vdd(vdd), .A(H_17_), .Y(_3965_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_3932_), .B(H_17_), .C(_3933_), .D(H_16_), .Y(_3966_) );
OAI21X1 OAI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .B(_3965_), .C(_3966_), .Y(_3967_) );
XOR2X1 XOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_19_), .Y(_3968_) );
INVX1 INVX1_501 ( .gnd(gnd), .vdd(vdd), .A(H_18_), .Y(_3969_) );
NAND2X1 NAND2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_3937_), .B(_3969_), .Y(_3970_) );
NAND2X1 NAND2X1_493 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_18_), .Y(_3971_) );
AOI21X1 AOI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_3970_), .B(_3971_), .C(_3968_), .Y(_3972_) );
NAND2X1 NAND2X1_494 ( .gnd(gnd), .vdd(vdd), .A(H_19_), .B(_3942_), .Y(_3894_) );
NAND2X1 NAND2X1_495 ( .gnd(gnd), .vdd(vdd), .A(H_18_), .B(_3937_), .Y(_3895_) );
OAI21X1 OAI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_3968_), .B(_3895_), .C(_3894_), .Y(_3896_) );
AOI21X1 AOI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_3967_), .B(_3972_), .C(_3896_), .Y(_3897_) );
INVX1 INVX1_502 ( .gnd(gnd), .vdd(vdd), .A(H_23_), .Y(_3898_) );
INVX1 INVX1_503 ( .gnd(gnd), .vdd(vdd), .A(H_22_), .Y(_3899_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3898_), .B(target[7]), .C(target[6]), .D(_3899_), .Y(_3900_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_3950_), .B(H_23_), .C(_3951_), .D(H_22_), .Y(_3901_) );
NOR2X1 NOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_3900_), .B(_3901_), .Y(_3902_) );
NAND2X1 NAND2X1_496 ( .gnd(gnd), .vdd(vdd), .A(H_21_), .B(_3957_), .Y(_3903_) );
NAND2X1 NAND2X1_497 ( .gnd(gnd), .vdd(vdd), .A(H_20_), .B(_3958_), .Y(_3904_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_3903_), .B(_3904_), .Y(_3905_) );
INVX1 INVX1_504 ( .gnd(gnd), .vdd(vdd), .A(H_20_), .Y(_3906_) );
NOR2X1 NOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(H_21_), .B(_3957_), .Y(_3907_) );
AOI21X1 AOI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_3906_), .C(_3907_), .Y(_3908_) );
NAND3X1 NAND3X1_937 ( .gnd(gnd), .vdd(vdd), .A(_3905_), .B(_3908_), .C(_3902_), .Y(_3909_) );
AOI21X1 AOI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_3903_), .B(_3904_), .C(_3907_), .Y(_3910_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3950_), .B(H_23_), .C(_3951_), .D(H_22_), .Y(_3911_) );
NOR2X1 NOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(H_23_), .B(_3950_), .Y(_3912_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3950_), .B(H_15_), .C(_3951_), .D(H_14_), .Y(_3913_) );
NOR2X1 NOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(H_15_), .B(_3950_), .Y(_3914_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3911_), .B(_3912_), .C(_3913_), .D(_3914_), .Y(_3915_) );
AOI21X1 AOI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_3902_), .B(_3910_), .C(_3915_), .Y(_3916_) );
OAI21X1 OAI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_3897_), .B(_3909_), .C(_3916_), .Y(_3917_) );
NOR2X1 NOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf0), .B(_3917__bF_buf2), .Y(_1_) );
INVX1 INVX1_505 ( .gnd(gnd), .vdd(vdd), .A(H_0_), .Y(_3918_) );
NOR3X1 NOR3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf2), .B(_3918_), .C(_3917__bF_buf1), .Y(_0__0_) );
INVX1 INVX1_506 ( .gnd(gnd), .vdd(vdd), .A(H_1_), .Y(_3919_) );
NOR3X1 NOR3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf2), .B(_3919_), .C(_3917__bF_buf0), .Y(_0__1_) );
INVX1 INVX1_507 ( .gnd(gnd), .vdd(vdd), .A(H_2_), .Y(_3920_) );
NOR3X1 NOR3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf3), .B(_3920_), .C(_3917__bF_buf4), .Y(_0__2_) );
INVX1 INVX1_508 ( .gnd(gnd), .vdd(vdd), .A(H_3_), .Y(_3921_) );
NOR3X1 NOR3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf4), .B(_3921_), .C(_3917__bF_buf0), .Y(_0__3_) );
INVX1 INVX1_509 ( .gnd(gnd), .vdd(vdd), .A(H_4_), .Y(_3922_) );
NOR3X1 NOR3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf3), .B(_3922_), .C(_3917__bF_buf4), .Y(_0__4_) );
INVX1 INVX1_510 ( .gnd(gnd), .vdd(vdd), .A(H_5_), .Y(_3923_) );
NOR3X1 NOR3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf2), .B(_3923_), .C(_3917__bF_buf0), .Y(_0__5_) );
INVX1 INVX1_511 ( .gnd(gnd), .vdd(vdd), .A(H_6_), .Y(_3924_) );
NOR3X1 NOR3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf3), .B(_3924_), .C(_3917__bF_buf4), .Y(_0__6_) );
INVX1 INVX1_512 ( .gnd(gnd), .vdd(vdd), .A(H_7_), .Y(_3925_) );
NOR3X1 NOR3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf3), .B(_3925_), .C(_3917__bF_buf4), .Y(_0__7_) );
INVX1 INVX1_513 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_3926_) );
NOR3X1 NOR3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf1), .B(_3926_), .C(_3917__bF_buf3), .Y(_0__8_) );
NOR3X1 NOR3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf3), .B(_3931_), .C(_3917__bF_buf4), .Y(_0__9_) );
NOR3X1 NOR3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf1), .B(_3938_), .C(_3917__bF_buf3), .Y(_0__10_) );
INVX1 INVX1_514 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_3927_) );
NOR3X1 NOR3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf1), .B(_3927_), .C(_3917__bF_buf3), .Y(_0__11_) );
NOR3X1 NOR3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf0), .B(_3955_), .C(_3917__bF_buf2), .Y(_0__12_) );
NOR3X1 NOR3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf4), .B(_3954_), .C(_3917__bF_buf1), .Y(_0__13_) );
NOR3X1 NOR3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf4), .B(_3948_), .C(_3917__bF_buf1), .Y(_0__14_) );
NOR3X1 NOR3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf4), .B(_3947_), .C(_3917__bF_buf0), .Y(_0__15_) );
INVX1 INVX1_515 ( .gnd(gnd), .vdd(vdd), .A(H_16_), .Y(_3928_) );
NOR3X1 NOR3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf2), .B(_3928_), .C(_3917__bF_buf0), .Y(_0__16_) );
NOR3X1 NOR3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf1), .B(_3965_), .C(_3917__bF_buf3), .Y(_0__17_) );
NOR3X1 NOR3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf1), .B(_3969_), .C(_3917__bF_buf3), .Y(_0__18_) );
INVX1 INVX1_516 ( .gnd(gnd), .vdd(vdd), .A(H_19_), .Y(_3929_) );
NOR3X1 NOR3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf2), .B(_3929_), .C(_3917__bF_buf1), .Y(_0__19_) );
NOR3X1 NOR3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf0), .B(_3906_), .C(_3917__bF_buf2), .Y(_0__20_) );
INVX1 INVX1_517 ( .gnd(gnd), .vdd(vdd), .A(H_21_), .Y(_3930_) );
NOR3X1 NOR3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf0), .B(_3930_), .C(_3917__bF_buf2), .Y(_0__21_) );
NOR3X1 NOR3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf0), .B(_3899_), .C(_3917__bF_buf2), .Y(_0__22_) );
NOR3X1 NOR3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_3964__bF_buf4), .B(_3898_), .C(_3917__bF_buf1), .Y(_0__23_) );
INVX1 INVX1_518 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[32]), .Y(_3973_) );
AOI21X1 AOI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(W_24_), .B(_3973_), .C(bloque_datos[80]), .Y(_3974_) );
OAI21X1 OAI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(W_24_), .B(_3973_), .C(_3974_), .Y(W_136_) );
INVX1 INVX1_519 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[33]), .Y(_3975_) );
AOI21X1 AOI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(W_25_), .B(_3975_), .C(bloque_datos[81]), .Y(_3976_) );
OAI21X1 OAI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(W_25_), .B(_3975_), .C(_3976_), .Y(W_137_) );
INVX1 INVX1_520 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[34]), .Y(_3977_) );
AOI21X1 AOI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(W_26_), .B(_3977_), .C(bloque_datos[82]), .Y(_3978_) );
OAI21X1 OAI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(W_26_), .B(_3977_), .C(_3978_), .Y(W_138_) );
INVX1 INVX1_521 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[35]), .Y(_3979_) );
AOI21X1 AOI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(W_27_), .B(_3979_), .C(bloque_datos[83]), .Y(_3980_) );
OAI21X1 OAI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(W_27_), .B(_3979_), .C(_3980_), .Y(W_139_) );
INVX1 INVX1_522 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[36]), .Y(_3981_) );
AOI21X1 AOI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(W_28_), .B(_3981_), .C(bloque_datos[84]), .Y(_3982_) );
OAI21X1 OAI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(W_28_), .B(_3981_), .C(_3982_), .Y(W_140_) );
INVX1 INVX1_523 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[37]), .Y(_3983_) );
AOI21X1 AOI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(W_29_), .B(_3983_), .C(bloque_datos[85]), .Y(_3984_) );
OAI21X1 OAI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(W_29_), .B(_3983_), .C(_3984_), .Y(W_141_) );
INVX1 INVX1_524 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[38]), .Y(_3985_) );
AOI21X1 AOI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(W_30_), .B(_3985_), .C(bloque_datos[86]), .Y(_3986_) );
OAI21X1 OAI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(W_30_), .B(_3985_), .C(_3986_), .Y(W_142_) );
INVX1 INVX1_525 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .Y(_3987_) );
AOI21X1 AOI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(W_31_), .B(_3987_), .C(bloque_datos[87]), .Y(_3988_) );
OAI21X1 OAI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(W_31_), .B(_3987_), .C(_3988_), .Y(W_143_) );
INVX1 INVX1_526 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[72]), .Y(_3989_) );
OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(W_16_), .B(bloque_datos[24]), .Y(_3990_) );
NAND2X1 NAND2X1_498 ( .gnd(gnd), .vdd(vdd), .A(W_16_), .B(bloque_datos[24]), .Y(_3991_) );
NAND2X1 NAND2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_3991_), .B(_3990_), .Y(_3992_) );
NAND2X1 NAND2X1_500 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .B(_3992_), .Y(W_128_) );
INVX1 INVX1_527 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[25]), .Y(_3993_) );
AOI21X1 AOI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(W_17_), .B(_3993_), .C(bloque_datos[73]), .Y(_3994_) );
OAI21X1 OAI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(W_17_), .B(_3993_), .C(_3994_), .Y(W_129_) );
INVX1 INVX1_528 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[74]), .Y(_3995_) );
OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(W_18_), .B(bloque_datos[26]), .Y(_3996_) );
NAND2X1 NAND2X1_501 ( .gnd(gnd), .vdd(vdd), .A(W_18_), .B(bloque_datos[26]), .Y(_3997_) );
NAND2X1 NAND2X1_502 ( .gnd(gnd), .vdd(vdd), .A(_3997_), .B(_3996_), .Y(_3998_) );
NAND2X1 NAND2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_3995_), .B(_3998_), .Y(W_130_) );
INVX1 INVX1_529 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[75]), .Y(_3999_) );
OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(W_19_), .B(bloque_datos[27]), .Y(_4000_) );
NAND2X1 NAND2X1_504 ( .gnd(gnd), .vdd(vdd), .A(W_19_), .B(bloque_datos[27]), .Y(_4001_) );
NAND2X1 NAND2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_4001_), .B(_4000_), .Y(_4002_) );
NAND2X1 NAND2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_3999_), .B(_4002_), .Y(W_131_) );
INVX2 INVX2_161 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[28]), .Y(_4003_) );
AOI21X1 AOI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(W_20_), .B(_4003_), .C(bloque_datos[76]), .Y(_4004_) );
OAI21X1 OAI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(W_20_), .B(_4003_), .C(_4004_), .Y(W_132_) );
INVX2 INVX2_162 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[29]), .Y(_4005_) );
AOI21X1 AOI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(W_21_), .B(_4005_), .C(bloque_datos[77]), .Y(_4006_) );
OAI21X1 OAI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(W_21_), .B(_4005_), .C(_4006_), .Y(W_133_) );
INVX2 INVX2_163 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[30]), .Y(_4007_) );
AOI21X1 AOI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(W_22_), .B(_4007_), .C(bloque_datos[78]), .Y(_4008_) );
OAI21X1 OAI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(W_22_), .B(_4007_), .C(_4008_), .Y(W_134_) );
INVX1 INVX1_530 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[31]), .Y(_4009_) );
AOI21X1 AOI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(W_23_), .B(_4009_), .C(bloque_datos[79]), .Y(_4010_) );
OAI21X1 OAI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(W_23_), .B(_4009_), .C(_4010_), .Y(W_135_) );
INVX1 INVX1_531 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(_4011_) );
INVX1 INVX1_532 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .Y(_4012_) );
OAI21X1 OAI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_4011_), .B(bloque_datos[40]), .C(_4012_), .Y(_4013_) );
AOI21X1 AOI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_4011_), .B(bloque_datos[40]), .C(_4013_), .Y(_4014_) );
INVX1 INVX1_533 ( .gnd(gnd), .vdd(vdd), .A(_4014_), .Y(W_144_) );
INVX1 INVX1_534 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(_4015_) );
INVX1 INVX1_535 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[89]), .Y(_4016_) );
OAI21X1 OAI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_4015_), .B(bloque_datos[41]), .C(_4016_), .Y(_4017_) );
AOI21X1 AOI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_4015_), .B(bloque_datos[41]), .C(_4017_), .Y(_4018_) );
INVX1 INVX1_536 ( .gnd(gnd), .vdd(vdd), .A(_4018_), .Y(W_145_) );
INVX1 INVX1_537 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[2]), .Y(_4019_) );
INVX1 INVX1_538 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[90]), .Y(_4020_) );
OAI21X1 OAI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_4019_), .B(bloque_datos[42]), .C(_4020_), .Y(_4021_) );
AOI21X1 AOI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_4019_), .B(bloque_datos[42]), .C(_4021_), .Y(_4022_) );
INVX1 INVX1_539 ( .gnd(gnd), .vdd(vdd), .A(_4022_), .Y(W_146_) );
INVX1 INVX1_540 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[3]), .Y(_4023_) );
INVX1 INVX1_541 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[91]), .Y(_4024_) );
OAI21X1 OAI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_4023_), .B(bloque_datos[43]), .C(_4024_), .Y(_4025_) );
AOI21X1 AOI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_4023_), .B(bloque_datos[43]), .C(_4025_), .Y(_4026_) );
INVX1 INVX1_542 ( .gnd(gnd), .vdd(vdd), .A(_4026_), .Y(W_147_) );
INVX1 INVX1_543 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[4]), .Y(_4027_) );
INVX1 INVX1_544 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[92]), .Y(_4028_) );
OAI21X1 OAI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_4027_), .B(bloque_datos[44]), .C(_4028_), .Y(_4029_) );
AOI21X1 AOI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_4027_), .B(bloque_datos[44]), .C(_4029_), .Y(_4030_) );
INVX1 INVX1_545 ( .gnd(gnd), .vdd(vdd), .A(_4030_), .Y(W_148_) );
INVX1 INVX1_546 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[5]), .Y(_4031_) );
INVX1 INVX1_547 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[93]), .Y(_4032_) );
OAI21X1 OAI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_4031_), .B(bloque_datos[45]), .C(_4032_), .Y(_4033_) );
AOI21X1 AOI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_4031_), .B(bloque_datos[45]), .C(_4033_), .Y(_4034_) );
INVX1 INVX1_548 ( .gnd(gnd), .vdd(vdd), .A(_4034_), .Y(W_149_) );
INVX1 INVX1_549 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[6]), .Y(_4035_) );
INVX1 INVX1_550 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[94]), .Y(_4036_) );
OAI21X1 OAI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(_4035_), .B(bloque_datos[46]), .C(_4036_), .Y(_4037_) );
AOI21X1 AOI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_4035_), .B(bloque_datos[46]), .C(_4037_), .Y(_4038_) );
INVX2 INVX2_164 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .Y(W_150_) );
INVX1 INVX1_551 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[7]), .Y(_4039_) );
INVX1 INVX1_552 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[95]), .Y(_4040_) );
OAI21X1 OAI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_4039_), .B(bloque_datos[47]), .C(_4040_), .Y(_4041_) );
AOI21X1 AOI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_4039_), .B(bloque_datos[47]), .C(_4041_), .Y(_4042_) );
INVX2 INVX2_165 ( .gnd(gnd), .vdd(vdd), .A(_4042_), .Y(W_151_) );
AOI21X1 AOI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_3991_), .B(_3990_), .C(bloque_datos[72]), .Y(_4043_) );
XNOR2X1 XNOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .B(bloque_datos[48]), .Y(_4044_) );
NAND2X1 NAND2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_4044_), .B(_4043_), .Y(W_152_) );
XOR2X1 XOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .B(bloque_datos[49]), .Y(_4045_) );
NOR2X1 NOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_4045_), .B(W_129_), .Y(_4046_) );
INVX1 INVX1_553 ( .gnd(gnd), .vdd(vdd), .A(_4046_), .Y(W_153_) );
AOI21X1 AOI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_3997_), .B(_3996_), .C(bloque_datos[74]), .Y(_4047_) );
XNOR2X1 XNOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .B(bloque_datos[50]), .Y(_4048_) );
NAND2X1 NAND2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_4048_), .B(_4047_), .Y(W_154_) );
AOI21X1 AOI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_4001_), .B(_4000_), .C(bloque_datos[75]), .Y(_4049_) );
XNOR2X1 XNOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .B(bloque_datos[51]), .Y(_4050_) );
NAND2X1 NAND2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_4050_), .B(_4049_), .Y(W_155_) );
INVX1 INVX1_554 ( .gnd(gnd), .vdd(vdd), .A(W_20_), .Y(_4051_) );
INVX1 INVX1_555 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[76]), .Y(_4052_) );
OAI21X1 OAI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_4051_), .B(bloque_datos[28]), .C(_4052_), .Y(_4053_) );
AOI21X1 AOI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_4051_), .B(bloque_datos[28]), .C(_4053_), .Y(_4054_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[12]), .B(bloque_datos[52]), .Y(_4055_) );
NOR2X1 NOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[12]), .B(bloque_datos[52]), .Y(_4056_) );
OAI21X1 OAI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_4055_), .B(_4056_), .C(_4054_), .Y(W_156_) );
XOR2X1 XOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[13]), .B(bloque_datos[53]), .Y(_4057_) );
NOR2X1 NOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_4057_), .B(W_133_), .Y(_4058_) );
INVX1 INVX1_556 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .Y(W_157_) );
XOR2X1 XOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[14]), .B(bloque_datos[54]), .Y(_4059_) );
NOR2X1 NOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_4059_), .B(W_134_), .Y(_4060_) );
INVX1 INVX1_557 ( .gnd(gnd), .vdd(vdd), .A(_4060_), .Y(W_158_) );
XOR2X1 XOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[15]), .B(bloque_datos[55]), .Y(_4061_) );
NOR2X1 NOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_4061_), .B(W_135_), .Y(_4062_) );
INVX1 INVX1_558 ( .gnd(gnd), .vdd(vdd), .A(_4062_), .Y(W_159_) );
XOR2X1 XOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(W_24_), .B(bloque_datos[32]), .Y(_4063_) );
NOR2X1 NOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .B(_4063_), .Y(_4064_) );
XNOR2X1 XNOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[16]), .B(bloque_datos[56]), .Y(_4065_) );
NAND2X1 NAND2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_4065_), .B(_4064_), .Y(W_160_) );
INVX1 INVX1_559 ( .gnd(gnd), .vdd(vdd), .A(W_25_), .Y(_4066_) );
INVX1 INVX1_560 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[81]), .Y(_4067_) );
OAI21X1 OAI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_4066_), .B(bloque_datos[33]), .C(_4067_), .Y(_4068_) );
AOI21X1 AOI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_4066_), .B(bloque_datos[33]), .C(_4068_), .Y(_4069_) );
XNOR2X1 XNOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .B(bloque_datos[57]), .Y(_4070_) );
NAND2X1 NAND2X1_511 ( .gnd(gnd), .vdd(vdd), .A(_4070_), .B(_4069_), .Y(W_161_) );
XOR2X1 XOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(W_26_), .B(bloque_datos[34]), .Y(_4071_) );
NOR2X1 NOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[82]), .B(_4071_), .Y(_4072_) );
XNOR2X1 XNOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .B(bloque_datos[58]), .Y(_4073_) );
NAND2X1 NAND2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_4073_), .B(_4072_), .Y(W_162_) );
XOR2X1 XOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(W_27_), .B(bloque_datos[35]), .Y(_4074_) );
NOR2X1 NOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[83]), .B(_4074_), .Y(_4075_) );
XNOR2X1 XNOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[19]), .B(bloque_datos[59]), .Y(_4076_) );
NAND2X1 NAND2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_4076_), .B(_4075_), .Y(W_163_) );
XOR2X1 XOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[20]), .B(bloque_datos[60]), .Y(_4077_) );
NOR2X1 NOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_4077_), .B(W_140_), .Y(_4078_) );
INVX1 INVX1_561 ( .gnd(gnd), .vdd(vdd), .A(_4078_), .Y(W_164_) );
XOR2X1 XOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[21]), .B(bloque_datos[61]), .Y(_4079_) );
NOR2X1 NOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_4079_), .B(W_141_), .Y(_4080_) );
INVX2 INVX2_166 ( .gnd(gnd), .vdd(vdd), .A(_4080_), .Y(W_165_) );
XOR2X1 XOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[22]), .B(bloque_datos[62]), .Y(_4081_) );
NOR2X1 NOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_4081_), .B(W_142_), .Y(_4082_) );
INVX2 INVX2_167 ( .gnd(gnd), .vdd(vdd), .A(_4082_), .Y(W_166_) );
XOR2X1 XOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[23]), .B(bloque_datos[63]), .Y(_4083_) );
NOR2X1 NOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_4083_), .B(W_143_), .Y(_4084_) );
INVX1 INVX1_562 ( .gnd(gnd), .vdd(vdd), .A(_4084_), .Y(W_167_) );
XNOR2X1 XNOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[24]), .B(bloque_datos[64]), .Y(_4085_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_4014_), .B(_4085_), .Y(_4086_) );
INVX2 INVX2_168 ( .gnd(gnd), .vdd(vdd), .A(_4086_), .Y(W_168_) );
XNOR2X1 XNOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[25]), .B(bloque_datos[65]), .Y(_4087_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_4018_), .B(_4087_), .Y(_4088_) );
INVX1 INVX1_563 ( .gnd(gnd), .vdd(vdd), .A(_4088_), .Y(W_169_) );
XNOR2X1 XNOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[26]), .B(bloque_datos[66]), .Y(_4089_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_4022_), .B(_4089_), .Y(_4090_) );
INVX1 INVX1_564 ( .gnd(gnd), .vdd(vdd), .A(_4090_), .Y(W_170_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[27]), .B(bloque_datos[67]), .Y(_4091_) );
NOR2X1 NOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[27]), .B(bloque_datos[67]), .Y(_4092_) );
OAI21X1 OAI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_4091_), .B(_4092_), .C(_4026_), .Y(W_171_) );
INVX2 INVX2_169 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[68]), .Y(_4093_) );
NOR2X1 NOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_4003_), .B(_4093_), .Y(_4094_) );
NOR2X1 NOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[28]), .B(bloque_datos[68]), .Y(_4095_) );
OAI21X1 OAI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_4094_), .B(_4095_), .C(_4030_), .Y(W_172_) );
INVX2 INVX2_170 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[69]), .Y(_4096_) );
NOR2X1 NOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_4005_), .B(_4096_), .Y(_4097_) );
NOR2X1 NOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[29]), .B(bloque_datos[69]), .Y(_4098_) );
OAI21X1 OAI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_4097_), .B(_4098_), .C(_4034_), .Y(W_173_) );
INVX2 INVX2_171 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[70]), .Y(_4099_) );
NOR2X1 NOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_4007_), .B(_4099_), .Y(_4100_) );
NOR2X1 NOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[30]), .B(bloque_datos[70]), .Y(_4101_) );
OAI21X1 OAI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_4100_), .B(_4101_), .C(_4038_), .Y(W_174_) );
XNOR2X1 XNOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[31]), .B(bloque_datos[71]), .Y(_4102_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_4042_), .B(_4102_), .Y(_4103_) );
INVX1 INVX1_565 ( .gnd(gnd), .vdd(vdd), .A(_4103_), .Y(W_175_) );
XNOR2X1 XNOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[32]), .B(bloque_datos[72]), .Y(_4104_) );
NAND3X1 NAND3X1_938 ( .gnd(gnd), .vdd(vdd), .A(_4044_), .B(_4104_), .C(_4043_), .Y(W_176_) );
INVX1 INVX1_566 ( .gnd(gnd), .vdd(vdd), .A(W_17_), .Y(_4105_) );
NAND2X1 NAND2X1_514 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[25]), .B(_4105_), .Y(_4106_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_3994_), .B(_4106_), .Y(_4107_) );
INVX1 INVX1_567 ( .gnd(gnd), .vdd(vdd), .A(_4045_), .Y(_4108_) );
XNOR2X1 XNOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[33]), .B(bloque_datos[73]), .Y(_4109_) );
NAND3X1 NAND3X1_939 ( .gnd(gnd), .vdd(vdd), .A(_4108_), .B(_4109_), .C(_4107_), .Y(W_177_) );
XNOR2X1 XNOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[34]), .B(bloque_datos[74]), .Y(_4110_) );
NAND3X1 NAND3X1_940 ( .gnd(gnd), .vdd(vdd), .A(_4048_), .B(_4110_), .C(_4047_), .Y(W_178_) );
XNOR2X1 XNOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[35]), .B(bloque_datos[75]), .Y(_4111_) );
NAND3X1 NAND3X1_941 ( .gnd(gnd), .vdd(vdd), .A(_4050_), .B(_4111_), .C(_4049_), .Y(W_179_) );
XOR2X1 XOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[36]), .B(bloque_datos[76]), .Y(_4112_) );
NOR2X1 NOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_4112_), .B(W_156_), .Y(_4113_) );
INVX1 INVX1_568 ( .gnd(gnd), .vdd(vdd), .A(_4113_), .Y(W_180_) );
INVX1 INVX1_569 ( .gnd(gnd), .vdd(vdd), .A(W_21_), .Y(_4114_) );
INVX1 INVX1_570 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[77]), .Y(_4115_) );
OAI21X1 OAI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_4114_), .B(bloque_datos[29]), .C(_4115_), .Y(_4116_) );
AOI21X1 AOI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_4114_), .B(bloque_datos[29]), .C(_4116_), .Y(_4117_) );
INVX1 INVX1_571 ( .gnd(gnd), .vdd(vdd), .A(_4057_), .Y(_4118_) );
XNOR2X1 XNOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[37]), .B(bloque_datos[77]), .Y(_4119_) );
NAND3X1 NAND3X1_942 ( .gnd(gnd), .vdd(vdd), .A(_4118_), .B(_4119_), .C(_4117_), .Y(W_181_) );
XNOR2X1 XNOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[38]), .B(bloque_datos[78]), .Y(_4120_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_4060_), .B(_4120_), .Y(_4121_) );
INVX2 INVX2_172 ( .gnd(gnd), .vdd(vdd), .A(_4121_), .Y(W_182_) );
XNOR2X1 XNOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .B(bloque_datos[79]), .Y(_4122_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_4062_), .B(_4122_), .Y(_4123_) );
INVX2 INVX2_173 ( .gnd(gnd), .vdd(vdd), .A(_4123_), .Y(W_183_) );
XNOR2X1 XNOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .B(bloque_datos[40]), .Y(_4124_) );
NAND3X1 NAND3X1_943 ( .gnd(gnd), .vdd(vdd), .A(_4065_), .B(_4124_), .C(_4064_), .Y(W_184_) );
XNOR2X1 XNOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[81]), .B(bloque_datos[41]), .Y(_4125_) );
NAND3X1 NAND3X1_944 ( .gnd(gnd), .vdd(vdd), .A(_4070_), .B(_4125_), .C(_4069_), .Y(W_185_) );
XNOR2X1 XNOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[82]), .B(bloque_datos[42]), .Y(_4126_) );
NAND3X1 NAND3X1_945 ( .gnd(gnd), .vdd(vdd), .A(_4073_), .B(_4126_), .C(_4072_), .Y(W_186_) );
XNOR2X1 XNOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[83]), .B(bloque_datos[43]), .Y(_4127_) );
NAND3X1 NAND3X1_946 ( .gnd(gnd), .vdd(vdd), .A(_4076_), .B(_4127_), .C(_4075_), .Y(W_187_) );
XNOR2X1 XNOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[84]), .B(bloque_datos[44]), .Y(_4128_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_4078_), .B(_4128_), .Y(_4129_) );
INVX1 INVX1_572 ( .gnd(gnd), .vdd(vdd), .A(_4129_), .Y(W_188_) );
XNOR2X1 XNOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[85]), .B(bloque_datos[45]), .Y(_4130_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_4080_), .B(_4130_), .Y(_4131_) );
INVX1 INVX1_573 ( .gnd(gnd), .vdd(vdd), .A(_4131_), .Y(W_189_) );
XNOR2X1 XNOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[86]), .B(bloque_datos[46]), .Y(_4132_) );
AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_4082_), .B(_4132_), .Y(_4133_) );
INVX1 INVX1_574 ( .gnd(gnd), .vdd(vdd), .A(_4133_), .Y(W_190_) );
XNOR2X1 XNOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[87]), .B(bloque_datos[47]), .Y(_4134_) );
AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_4084_), .B(_4134_), .Y(_4135_) );
INVX1 INVX1_575 ( .gnd(gnd), .vdd(vdd), .A(_4135_), .Y(W_191_) );
AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .B(bloque_datos[48]), .Y(_4136_) );
NOR2X1 NOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .B(bloque_datos[48]), .Y(_4137_) );
OAI21X1 OAI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_4136_), .B(_4137_), .C(_4086_), .Y(W_192_) );
AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[89]), .B(bloque_datos[49]), .Y(_4138_) );
NOR2X1 NOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[89]), .B(bloque_datos[49]), .Y(_4139_) );
OAI21X1 OAI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_4138_), .B(_4139_), .C(_4088_), .Y(W_193_) );
AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[90]), .B(bloque_datos[50]), .Y(_4140_) );
NOR2X1 NOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[90]), .B(bloque_datos[50]), .Y(_4141_) );
OAI21X1 OAI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_4140_), .B(_4141_), .C(_4090_), .Y(W_194_) );
OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(W_171_), .B(bloque_datos[51]), .Y(W_195_) );
NOR2X1 NOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[52]), .B(W_172_), .Y(_4142_) );
INVX1 INVX1_576 ( .gnd(gnd), .vdd(vdd), .A(_4142_), .Y(W_196_) );
NOR2X1 NOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[53]), .B(W_173_), .Y(_4143_) );
INVX1 INVX1_577 ( .gnd(gnd), .vdd(vdd), .A(_4143_), .Y(W_197_) );
OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(W_174_), .B(bloque_datos[54]), .Y(W_198_) );
XNOR2X1 XNOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[95]), .B(bloque_datos[55]), .Y(_4144_) );
NAND2X1 NAND2X1_515 ( .gnd(gnd), .vdd(vdd), .A(_4144_), .B(_4103_), .Y(W_199_) );
NAND2X1 NAND2X1_516 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[56]), .B(W_128_), .Y(_4145_) );
INVX1 INVX1_578 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[56]), .Y(_4146_) );
NAND2X1 NAND2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_4146_), .B(_4043_), .Y(_4147_) );
AOI21X1 AOI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_4147_), .B(_4145_), .C(W_176_), .Y(_4148_) );
INVX2 INVX2_174 ( .gnd(gnd), .vdd(vdd), .A(_4148_), .Y(W_200_) );
NAND2X1 NAND2X1_518 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[57]), .B(W_129_), .Y(_4149_) );
OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(W_129_), .B(bloque_datos[57]), .Y(_4150_) );
AOI21X1 AOI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_4149_), .B(_4150_), .C(W_177_), .Y(_4151_) );
INVX1 INVX1_579 ( .gnd(gnd), .vdd(vdd), .A(_4151_), .Y(W_201_) );
NAND2X1 NAND2X1_519 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[58]), .B(W_130_), .Y(_4152_) );
INVX1 INVX1_580 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[58]), .Y(_4153_) );
NAND2X1 NAND2X1_520 ( .gnd(gnd), .vdd(vdd), .A(_4153_), .B(_4047_), .Y(_4154_) );
AOI21X1 AOI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_4154_), .B(_4152_), .C(W_178_), .Y(_4155_) );
INVX1 INVX1_581 ( .gnd(gnd), .vdd(vdd), .A(_4155_), .Y(W_202_) );
NAND2X1 NAND2X1_521 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[59]), .B(W_131_), .Y(_4156_) );
INVX1 INVX1_582 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[59]), .Y(_4157_) );
NAND2X1 NAND2X1_522 ( .gnd(gnd), .vdd(vdd), .A(_4157_), .B(_4049_), .Y(_4158_) );
AOI21X1 AOI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_4158_), .B(_4156_), .C(W_179_), .Y(_4159_) );
INVX1 INVX1_583 ( .gnd(gnd), .vdd(vdd), .A(_4159_), .Y(W_203_) );
XNOR2X1 XNOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(W_132_), .B(bloque_datos[60]), .Y(_4160_) );
NAND2X1 NAND2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_4160_), .B(_4113_), .Y(W_204_) );
NAND2X1 NAND2X1_524 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[61]), .B(W_133_), .Y(_4161_) );
OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(W_133_), .B(bloque_datos[61]), .Y(_4162_) );
AOI21X1 AOI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_4161_), .B(_4162_), .C(W_181_), .Y(_4163_) );
INVX1 INVX1_584 ( .gnd(gnd), .vdd(vdd), .A(_4163_), .Y(W_205_) );
INVX2 INVX2_175 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[62]), .Y(_4164_) );
NAND2X1 NAND2X1_525 ( .gnd(gnd), .vdd(vdd), .A(_4164_), .B(_4121_), .Y(W_206_) );
INVX2 INVX2_176 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[63]), .Y(_4165_) );
NAND2X1 NAND2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_4165_), .B(_4123_), .Y(W_207_) );
OAI21X1 OAI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_4063_), .B(bloque_datos[80]), .C(bloque_datos[64]), .Y(_4166_) );
OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(W_136_), .B(bloque_datos[64]), .Y(_4167_) );
AOI21X1 AOI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_4166_), .B(_4167_), .C(W_184_), .Y(_4168_) );
INVX2 INVX2_177 ( .gnd(gnd), .vdd(vdd), .A(_4168_), .Y(W_208_) );
NAND2X1 NAND2X1_527 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[65]), .B(W_137_), .Y(_4169_) );
OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(W_137_), .B(bloque_datos[65]), .Y(_4170_) );
AOI21X1 AOI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_4169_), .B(_4170_), .C(W_185_), .Y(_4171_) );
INVX1 INVX1_585 ( .gnd(gnd), .vdd(vdd), .A(_4171_), .Y(W_209_) );
OAI21X1 OAI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_4071_), .B(bloque_datos[82]), .C(bloque_datos[66]), .Y(_4172_) );
OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(W_138_), .B(bloque_datos[66]), .Y(_4173_) );
AOI21X1 AOI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_4172_), .B(_4173_), .C(W_186_), .Y(_4174_) );
INVX1 INVX1_586 ( .gnd(gnd), .vdd(vdd), .A(_4174_), .Y(W_210_) );
OAI21X1 OAI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(_4074_), .B(bloque_datos[83]), .C(bloque_datos[67]), .Y(_4175_) );
OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(W_139_), .B(bloque_datos[67]), .Y(_4176_) );
AOI21X1 AOI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_4175_), .B(_4176_), .C(W_187_), .Y(_4177_) );
INVX2 INVX2_178 ( .gnd(gnd), .vdd(vdd), .A(_4177_), .Y(W_211_) );
NAND2X1 NAND2X1_528 ( .gnd(gnd), .vdd(vdd), .A(_4093_), .B(_4129_), .Y(W_212_) );
NAND2X1 NAND2X1_529 ( .gnd(gnd), .vdd(vdd), .A(_4096_), .B(_4131_), .Y(W_213_) );
NAND2X1 NAND2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_4099_), .B(_4133_), .Y(W_214_) );
INVX1 INVX1_587 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[71]), .Y(_4178_) );
NAND2X1 NAND2X1_531 ( .gnd(gnd), .vdd(vdd), .A(_4178_), .B(_4135_), .Y(W_215_) );
OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(W_192_), .B(bloque_datos[72]), .Y(W_216_) );
OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(W_193_), .B(bloque_datos[73]), .Y(W_217_) );
OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(W_194_), .B(bloque_datos[74]), .Y(W_218_) );
OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(W_195_), .B(bloque_datos[75]), .Y(W_219_) );
NAND2X1 NAND2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_4052_), .B(_4142_), .Y(W_220_) );
NAND2X1 NAND2X1_533 ( .gnd(gnd), .vdd(vdd), .A(_4115_), .B(_4143_), .Y(W_221_) );
OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(W_198_), .B(bloque_datos[78]), .Y(W_222_) );
OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(W_199_), .B(bloque_datos[79]), .Y(W_223_) );
XNOR2X1 XNOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(W_152_), .B(bloque_datos[80]), .Y(_4179_) );
NAND2X1 NAND2X1_534 ( .gnd(gnd), .vdd(vdd), .A(_4148_), .B(_4179_), .Y(W_224_) );
OAI21X1 OAI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(W_129_), .B(_4045_), .C(bloque_datos[81]), .Y(_4180_) );
NAND3X1 NAND3X1_947 ( .gnd(gnd), .vdd(vdd), .A(_4067_), .B(_4108_), .C(_4107_), .Y(_4181_) );
NAND2X1 NAND2X1_535 ( .gnd(gnd), .vdd(vdd), .A(_4180_), .B(_4181_), .Y(_4182_) );
NAND2X1 NAND2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_4182_), .B(_4151_), .Y(W_225_) );
XNOR2X1 XNOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(W_154_), .B(bloque_datos[82]), .Y(_4183_) );
NAND2X1 NAND2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_4155_), .B(_4183_), .Y(W_226_) );
XNOR2X1 XNOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(W_155_), .B(bloque_datos[83]), .Y(_4184_) );
NAND2X1 NAND2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_4159_), .B(_4184_), .Y(W_227_) );
INVX1 INVX1_588 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[84]), .Y(_4185_) );
NAND3X1 NAND3X1_948 ( .gnd(gnd), .vdd(vdd), .A(_4185_), .B(_4160_), .C(_4113_), .Y(W_228_) );
OAI21X1 OAI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(W_133_), .B(_4057_), .C(bloque_datos[85]), .Y(_4186_) );
INVX1 INVX1_589 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[85]), .Y(_4187_) );
NAND3X1 NAND3X1_949 ( .gnd(gnd), .vdd(vdd), .A(_4187_), .B(_4118_), .C(_4117_), .Y(_4188_) );
NAND2X1 NAND2X1_539 ( .gnd(gnd), .vdd(vdd), .A(_4186_), .B(_4188_), .Y(_4189_) );
NAND2X1 NAND2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_4189_), .B(_4163_), .Y(W_229_) );
INVX1 INVX1_590 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[86]), .Y(_4190_) );
NAND3X1 NAND3X1_950 ( .gnd(gnd), .vdd(vdd), .A(_4190_), .B(_4164_), .C(_4121_), .Y(W_230_) );
INVX1 INVX1_591 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[87]), .Y(_4191_) );
NAND3X1 NAND3X1_951 ( .gnd(gnd), .vdd(vdd), .A(_4191_), .B(_4165_), .C(_4123_), .Y(W_231_) );
AOI21X1 AOI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_4065_), .B(_4064_), .C(_4012_), .Y(_4192_) );
NOR2X1 NOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .B(W_160_), .Y(_4193_) );
OAI21X1 OAI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_4193_), .B(_4192_), .C(_4168_), .Y(W_232_) );
AOI21X1 AOI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_4070_), .B(_4069_), .C(_4016_), .Y(_4194_) );
NOR2X1 NOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[89]), .B(W_161_), .Y(_4195_) );
OAI21X1 OAI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_4194_), .B(_4195_), .C(_4171_), .Y(W_233_) );
AOI21X1 AOI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_4073_), .B(_4072_), .C(_4020_), .Y(_4196_) );
NOR2X1 NOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[90]), .B(W_162_), .Y(_4197_) );
OAI21X1 OAI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_4197_), .B(_4196_), .C(_4174_), .Y(W_234_) );
AOI21X1 AOI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_4076_), .B(_4075_), .C(_4024_), .Y(_4198_) );
NOR2X1 NOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[91]), .B(W_163_), .Y(_4199_) );
OAI21X1 OAI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_4199_), .B(_4198_), .C(_4177_), .Y(W_235_) );
NAND3X1 NAND3X1_952 ( .gnd(gnd), .vdd(vdd), .A(_4028_), .B(_4093_), .C(_4129_), .Y(W_236_) );
NAND3X1 NAND3X1_953 ( .gnd(gnd), .vdd(vdd), .A(_4032_), .B(_4096_), .C(_4131_), .Y(W_237_) );
NAND3X1 NAND3X1_954 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .B(_4099_), .C(_4133_), .Y(W_238_) );
NAND3X1 NAND3X1_955 ( .gnd(gnd), .vdd(vdd), .A(_4040_), .B(_4178_), .C(_4135_), .Y(W_239_) );
OR2X2 OR2X2_90 ( .gnd(gnd), .vdd(vdd), .A(W_192_), .B(W_128_), .Y(W_240_) );
OR2X2 OR2X2_91 ( .gnd(gnd), .vdd(vdd), .A(W_193_), .B(W_129_), .Y(W_241_) );
OR2X2 OR2X2_92 ( .gnd(gnd), .vdd(vdd), .A(W_194_), .B(W_130_), .Y(W_242_) );
OR2X2 OR2X2_93 ( .gnd(gnd), .vdd(vdd), .A(W_195_), .B(W_131_), .Y(W_243_) );
NAND2X1 NAND2X1_541 ( .gnd(gnd), .vdd(vdd), .A(_4054_), .B(_4142_), .Y(W_244_) );
NAND2X1 NAND2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_4117_), .B(_4143_), .Y(W_245_) );
OR2X2 OR2X2_94 ( .gnd(gnd), .vdd(vdd), .A(W_198_), .B(W_134_), .Y(W_246_) );
OR2X2 OR2X2_95 ( .gnd(gnd), .vdd(vdd), .A(W_199_), .B(W_135_), .Y(W_247_) );
XNOR2X1 XNOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(W_176_), .B(W_136_), .Y(_4200_) );
NAND3X1 NAND3X1_956 ( .gnd(gnd), .vdd(vdd), .A(_4148_), .B(_4179_), .C(_4200_), .Y(W_248_) );
NAND3X1 NAND3X1_957 ( .gnd(gnd), .vdd(vdd), .A(_4069_), .B(_4182_), .C(_4151_), .Y(W_249_) );
XNOR2X1 XNOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(W_178_), .B(W_138_), .Y(_4201_) );
NAND3X1 NAND3X1_958 ( .gnd(gnd), .vdd(vdd), .A(_4155_), .B(_4183_), .C(_4201_), .Y(W_250_) );
XNOR2X1 XNOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(W_179_), .B(W_139_), .Y(_4202_) );
NAND3X1 NAND3X1_959 ( .gnd(gnd), .vdd(vdd), .A(_4159_), .B(_4184_), .C(_4202_), .Y(W_251_) );
INVX1 INVX1_592 ( .gnd(gnd), .vdd(vdd), .A(W_140_), .Y(_4203_) );
NAND3X1 NAND3X1_960 ( .gnd(gnd), .vdd(vdd), .A(_4203_), .B(_4160_), .C(_4113_), .Y(W_252_) );
INVX1 INVX1_593 ( .gnd(gnd), .vdd(vdd), .A(W_141_), .Y(_4204_) );
NAND3X1 NAND3X1_961 ( .gnd(gnd), .vdd(vdd), .A(_4204_), .B(_4189_), .C(_4163_), .Y(W_253_) );
INVX1 INVX1_594 ( .gnd(gnd), .vdd(vdd), .A(W_142_), .Y(_4205_) );
NAND3X1 NAND3X1_962 ( .gnd(gnd), .vdd(vdd), .A(_4164_), .B(_4205_), .C(_4121_), .Y(W_254_) );
INVX1 INVX1_595 ( .gnd(gnd), .vdd(vdd), .A(W_143_), .Y(_4206_) );
NAND3X1 NAND3X1_963 ( .gnd(gnd), .vdd(vdd), .A(_4165_), .B(_4206_), .C(_4123_), .Y(W_255_) );
BUFX2 BUFX2_126 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__24_) );
BUFX2 BUFX2_127 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__25_) );
BUFX2 BUFX2_128 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__26_) );
BUFX2 BUFX2_129 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__27_) );
BUFX2 BUFX2_130 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__28_) );
BUFX2 BUFX2_131 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__29_) );
BUFX2 BUFX2_132 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__30_) );
BUFX2 BUFX2_133 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__31_) );
BUFX2 BUFX2_134 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__32_) );
BUFX2 BUFX2_135 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__33_) );
BUFX2 BUFX2_136 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__34_) );
BUFX2 BUFX2_137 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__35_) );
BUFX2 BUFX2_138 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__36_) );
BUFX2 BUFX2_139 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__37_) );
BUFX2 BUFX2_140 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__38_) );
BUFX2 BUFX2_141 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__39_) );
BUFX2 BUFX2_142 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__40_) );
BUFX2 BUFX2_143 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__41_) );
BUFX2 BUFX2_144 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__42_) );
BUFX2 BUFX2_145 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__43_) );
BUFX2 BUFX2_146 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__44_) );
BUFX2 BUFX2_147 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__45_) );
BUFX2 BUFX2_148 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__46_) );
BUFX2 BUFX2_149 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__47_) );
BUFX2 BUFX2_150 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__48_) );
BUFX2 BUFX2_151 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__49_) );
BUFX2 BUFX2_152 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__50_) );
BUFX2 BUFX2_153 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__51_) );
BUFX2 BUFX2_154 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__52_) );
BUFX2 BUFX2_155 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__53_) );
BUFX2 BUFX2_156 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__54_) );
BUFX2 BUFX2_157 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__55_) );
BUFX2 BUFX2_158 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__56_) );
BUFX2 BUFX2_159 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__57_) );
BUFX2 BUFX2_160 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__58_) );
BUFX2 BUFX2_161 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__59_) );
BUFX2 BUFX2_162 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__60_) );
BUFX2 BUFX2_163 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__61_) );
BUFX2 BUFX2_164 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__62_) );
BUFX2 BUFX2_165 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__63_) );
BUFX2 BUFX2_166 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__64_) );
BUFX2 BUFX2_167 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__65_) );
BUFX2 BUFX2_168 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__66_) );
BUFX2 BUFX2_169 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__67_) );
BUFX2 BUFX2_170 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__68_) );
BUFX2 BUFX2_171 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__69_) );
BUFX2 BUFX2_172 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__70_) );
BUFX2 BUFX2_173 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__71_) );
BUFX2 BUFX2_174 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__72_) );
BUFX2 BUFX2_175 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__73_) );
BUFX2 BUFX2_176 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__74_) );
BUFX2 BUFX2_177 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__75_) );
BUFX2 BUFX2_178 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__76_) );
BUFX2 BUFX2_179 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__77_) );
BUFX2 BUFX2_180 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__78_) );
BUFX2 BUFX2_181 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__79_) );
BUFX2 BUFX2_182 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__80_) );
BUFX2 BUFX2_183 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__81_) );
BUFX2 BUFX2_184 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__82_) );
BUFX2 BUFX2_185 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__83_) );
BUFX2 BUFX2_186 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__84_) );
BUFX2 BUFX2_187 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__85_) );
BUFX2 BUFX2_188 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__86_) );
BUFX2 BUFX2_189 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__87_) );
BUFX2 BUFX2_190 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__88_) );
BUFX2 BUFX2_191 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__89_) );
BUFX2 BUFX2_192 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__90_) );
BUFX2 BUFX2_193 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__91_) );
BUFX2 BUFX2_194 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__92_) );
BUFX2 BUFX2_195 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__93_) );
BUFX2 BUFX2_196 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__94_) );
BUFX2 BUFX2_197 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__95_) );
BUFX2 BUFX2_198 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__96_) );
BUFX2 BUFX2_199 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__97_) );
BUFX2 BUFX2_200 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__98_) );
BUFX2 BUFX2_201 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__99_) );
BUFX2 BUFX2_202 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__100_) );
BUFX2 BUFX2_203 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__101_) );
BUFX2 BUFX2_204 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__102_) );
BUFX2 BUFX2_205 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__103_) );
BUFX2 BUFX2_206 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__104_) );
BUFX2 BUFX2_207 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__105_) );
BUFX2 BUFX2_208 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__106_) );
BUFX2 BUFX2_209 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__107_) );
BUFX2 BUFX2_210 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__108_) );
BUFX2 BUFX2_211 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__109_) );
BUFX2 BUFX2_212 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__110_) );
BUFX2 BUFX2_213 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__111_) );
BUFX2 BUFX2_214 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__112_) );
BUFX2 BUFX2_215 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__113_) );
BUFX2 BUFX2_216 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__114_) );
BUFX2 BUFX2_217 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__115_) );
BUFX2 BUFX2_218 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__116_) );
BUFX2 BUFX2_219 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__117_) );
BUFX2 BUFX2_220 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__118_) );
BUFX2 BUFX2_221 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__119_) );
BUFX2 BUFX2_222 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__120_) );
BUFX2 BUFX2_223 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__121_) );
BUFX2 BUFX2_224 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__122_) );
BUFX2 BUFX2_225 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_0__123_) );
BUFX2 BUFX2_226 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(H_8_) );
BUFX2 BUFX2_227 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(H_9_) );
BUFX2 BUFX2_228 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(H_10_) );
BUFX2 BUFX2_229 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(H_11_) );
BUFX2 BUFX2_230 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(W_32_) );
BUFX2 BUFX2_231 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(W_33_) );
BUFX2 BUFX2_232 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[2]), .Y(W_34_) );
BUFX2 BUFX2_233 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[3]), .Y(W_35_) );
BUFX2 BUFX2_234 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[4]), .Y(W_36_) );
BUFX2 BUFX2_235 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[5]), .Y(W_37_) );
BUFX2 BUFX2_236 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[6]), .Y(W_38_) );
BUFX2 BUFX2_237 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[7]), .Y(W_39_) );
BUFX2 BUFX2_238 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .Y(W_40_) );
BUFX2 BUFX2_239 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .Y(W_41_) );
BUFX2 BUFX2_240 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .Y(W_42_) );
BUFX2 BUFX2_241 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .Y(W_43_) );
BUFX2 BUFX2_242 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[12]), .Y(W_44_) );
BUFX2 BUFX2_243 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[13]), .Y(W_45_) );
BUFX2 BUFX2_244 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[14]), .Y(W_46_) );
BUFX2 BUFX2_245 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[15]), .Y(W_47_) );
BUFX2 BUFX2_246 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[16]), .Y(W_48_) );
BUFX2 BUFX2_247 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .Y(W_49_) );
BUFX2 BUFX2_248 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .Y(W_50_) );
BUFX2 BUFX2_249 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[19]), .Y(W_51_) );
BUFX2 BUFX2_250 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[20]), .Y(W_52_) );
BUFX2 BUFX2_251 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[21]), .Y(W_53_) );
BUFX2 BUFX2_252 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[22]), .Y(W_54_) );
BUFX2 BUFX2_253 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[23]), .Y(W_55_) );
BUFX2 BUFX2_254 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[24]), .Y(W_56_) );
BUFX2 BUFX2_255 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[25]), .Y(W_57_) );
BUFX2 BUFX2_256 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[26]), .Y(W_58_) );
BUFX2 BUFX2_257 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[27]), .Y(W_59_) );
BUFX2 BUFX2_258 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[28]), .Y(W_60_) );
BUFX2 BUFX2_259 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[29]), .Y(W_61_) );
BUFX2 BUFX2_260 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[30]), .Y(W_62_) );
BUFX2 BUFX2_261 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[31]), .Y(W_63_) );
BUFX2 BUFX2_262 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[32]), .Y(W_64_) );
BUFX2 BUFX2_263 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[33]), .Y(W_65_) );
BUFX2 BUFX2_264 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[34]), .Y(W_66_) );
BUFX2 BUFX2_265 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[35]), .Y(W_67_) );
BUFX2 BUFX2_266 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[36]), .Y(W_68_) );
BUFX2 BUFX2_267 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[37]), .Y(W_69_) );
BUFX2 BUFX2_268 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[38]), .Y(W_70_) );
BUFX2 BUFX2_269 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .Y(W_71_) );
BUFX2 BUFX2_270 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[40]), .Y(W_72_) );
BUFX2 BUFX2_271 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[41]), .Y(W_73_) );
BUFX2 BUFX2_272 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[42]), .Y(W_74_) );
BUFX2 BUFX2_273 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[43]), .Y(W_75_) );
BUFX2 BUFX2_274 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[44]), .Y(W_76_) );
BUFX2 BUFX2_275 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[45]), .Y(W_77_) );
BUFX2 BUFX2_276 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[46]), .Y(W_78_) );
BUFX2 BUFX2_277 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[47]), .Y(W_79_) );
BUFX2 BUFX2_278 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[48]), .Y(W_80_) );
BUFX2 BUFX2_279 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[49]), .Y(W_81_) );
BUFX2 BUFX2_280 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[50]), .Y(W_82_) );
BUFX2 BUFX2_281 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[51]), .Y(W_83_) );
BUFX2 BUFX2_282 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[52]), .Y(W_84_) );
BUFX2 BUFX2_283 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[53]), .Y(W_85_) );
BUFX2 BUFX2_284 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[54]), .Y(W_86_) );
BUFX2 BUFX2_285 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[55]), .Y(W_87_) );
BUFX2 BUFX2_286 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[56]), .Y(W_88_) );
BUFX2 BUFX2_287 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[57]), .Y(W_89_) );
BUFX2 BUFX2_288 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[58]), .Y(W_90_) );
BUFX2 BUFX2_289 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[59]), .Y(W_91_) );
BUFX2 BUFX2_290 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[60]), .Y(W_92_) );
BUFX2 BUFX2_291 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[61]), .Y(W_93_) );
BUFX2 BUFX2_292 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[62]), .Y(W_94_) );
BUFX2 BUFX2_293 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[63]), .Y(W_95_) );
BUFX2 BUFX2_294 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[64]), .Y(W_96_) );
BUFX2 BUFX2_295 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[65]), .Y(W_97_) );
BUFX2 BUFX2_296 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[66]), .Y(W_98_) );
BUFX2 BUFX2_297 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[67]), .Y(W_99_) );
BUFX2 BUFX2_298 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[68]), .Y(W_100_) );
BUFX2 BUFX2_299 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[69]), .Y(W_101_) );
BUFX2 BUFX2_300 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[70]), .Y(W_102_) );
BUFX2 BUFX2_301 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[71]), .Y(W_103_) );
BUFX2 BUFX2_302 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[72]), .Y(W_104_) );
BUFX2 BUFX2_303 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[73]), .Y(W_105_) );
BUFX2 BUFX2_304 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[74]), .Y(W_106_) );
BUFX2 BUFX2_305 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[75]), .Y(W_107_) );
BUFX2 BUFX2_306 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[76]), .Y(W_108_) );
BUFX2 BUFX2_307 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[77]), .Y(W_109_) );
BUFX2 BUFX2_308 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[78]), .Y(W_110_) );
BUFX2 BUFX2_309 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[79]), .Y(W_111_) );
BUFX2 BUFX2_310 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .Y(W_112_) );
BUFX2 BUFX2_311 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[81]), .Y(W_113_) );
BUFX2 BUFX2_312 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[82]), .Y(W_114_) );
BUFX2 BUFX2_313 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[83]), .Y(W_115_) );
BUFX2 BUFX2_314 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[84]), .Y(W_116_) );
BUFX2 BUFX2_315 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[85]), .Y(W_117_) );
BUFX2 BUFX2_316 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[86]), .Y(W_118_) );
BUFX2 BUFX2_317 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[87]), .Y(W_119_) );
BUFX2 BUFX2_318 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .Y(W_120_) );
BUFX2 BUFX2_319 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[89]), .Y(W_121_) );
BUFX2 BUFX2_320 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[90]), .Y(W_122_) );
BUFX2 BUFX2_321 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[91]), .Y(W_123_) );
BUFX2 BUFX2_322 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[92]), .Y(W_124_) );
BUFX2 BUFX2_323 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[93]), .Y(W_125_) );
BUFX2 BUFX2_324 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[94]), .Y(W_126_) );
BUFX2 BUFX2_325 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[95]), .Y(W_127_) );
endmodule
