module micro_ucr_hash_mod ( gnd, vdd, clk, bloque_datos, inicio, nonce_iniciales, target, bounty_out, terminado_out);

input gnd, vdd;
input clk;
input inicio;
output terminado_out;
input [95:0] bloque_datos;
input [127:0] nonce_iniciales;
input [7:0] target;
output [23:0] bounty_out;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[83]), .Y(bloque_datos_83_bF_buf5_) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[83]), .Y(bloque_datos_83_bF_buf4_) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[83]), .Y(bloque_datos_83_bF_buf3_) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[83]), .Y(bloque_datos_83_bF_buf2_) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[83]), .Y(bloque_datos_83_bF_buf1_) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[83]), .Y(bloque_datos_83_bF_buf0_) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(_12797_), .Y(_12797__bF_buf4) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(_12797_), .Y(_12797__bF_buf3) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(_12797_), .Y(_12797__bF_buf2) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(_12797_), .Y(_12797__bF_buf1) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(_12797_), .Y(_12797__bF_buf0) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[42]), .Y(bloque_datos_42_bF_buf3_) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[42]), .Y(bloque_datos_42_bF_buf2_) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[42]), .Y(bloque_datos_42_bF_buf1_) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[42]), .Y(bloque_datos_42_bF_buf0_) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .Y(bloque_datos_80_bF_buf5_) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .Y(bloque_datos_80_bF_buf4_) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .Y(bloque_datos_80_bF_buf3_) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .Y(bloque_datos_80_bF_buf2_) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .Y(bloque_datos_80_bF_buf1_) );
BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[80]), .Y(bloque_datos_80_bF_buf0_) );
BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[77]), .Y(bloque_datos_77_bF_buf4_) );
BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[77]), .Y(bloque_datos_77_bF_buf3_) );
BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[77]), .Y(bloque_datos_77_bF_buf2_) );
BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[77]), .Y(bloque_datos_77_bF_buf1_) );
BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[77]), .Y(bloque_datos_77_bF_buf0_) );
BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(_16933_), .Y(_16933__bF_buf3) );
BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(_16933_), .Y(_16933__bF_buf2) );
BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(_16933_), .Y(_16933__bF_buf1) );
BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(_16933_), .Y(_16933__bF_buf0) );
BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado), .Y(module_1_comparador_target_hash_0_terminado_bF_buf6) );
BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado), .Y(module_1_comparador_target_hash_0_terminado_bF_buf5) );
BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado), .Y(module_1_comparador_target_hash_0_terminado_bF_buf4) );
BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado), .Y(module_1_comparador_target_hash_0_terminado_bF_buf3) );
BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado), .Y(module_1_comparador_target_hash_0_terminado_bF_buf2) );
BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado), .Y(module_1_comparador_target_hash_0_terminado_bF_buf1) );
BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado), .Y(module_1_comparador_target_hash_0_terminado_bF_buf0) );
BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[36]), .Y(bloque_datos_36_bF_buf3_) );
BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[36]), .Y(bloque_datos_36_bF_buf2_) );
BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[36]), .Y(bloque_datos_36_bF_buf1_) );
BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[36]), .Y(bloque_datos_36_bF_buf0_) );
BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado), .Y(module_3_comparador_target_hash_0_terminado_bF_buf6) );
BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado), .Y(module_3_comparador_target_hash_0_terminado_bF_buf5) );
BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado), .Y(module_3_comparador_target_hash_0_terminado_bF_buf4) );
BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado), .Y(module_3_comparador_target_hash_0_terminado_bF_buf3) );
BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado), .Y(module_3_comparador_target_hash_0_terminado_bF_buf2) );
BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado), .Y(module_3_comparador_target_hash_0_terminado_bF_buf1) );
BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado), .Y(module_3_comparador_target_hash_0_terminado_bF_buf0) );
BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[74]), .Y(bloque_datos_74_bF_buf4_) );
BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[74]), .Y(bloque_datos_74_bF_buf3_) );
BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[74]), .Y(bloque_datos_74_bF_buf2_) );
BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[74]), .Y(bloque_datos_74_bF_buf1_) );
BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[74]), .Y(bloque_datos_74_bF_buf0_) );
BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[33]), .Y(bloque_datos_33_bF_buf3_) );
BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[33]), .Y(bloque_datos_33_bF_buf2_) );
BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[33]), .Y(bloque_datos_33_bF_buf1_) );
BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[33]), .Y(bloque_datos_33_bF_buf0_) );
BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[71]), .Y(bloque_datos_71_bF_buf3_) );
BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[71]), .Y(bloque_datos_71_bF_buf2_) );
BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[71]), .Y(bloque_datos_71_bF_buf1_) );
BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[71]), .Y(bloque_datos_71_bF_buf0_) );
BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[6]), .Y(bloque_datos_6_bF_buf3_) );
BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[6]), .Y(bloque_datos_6_bF_buf2_) );
BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[6]), .Y(bloque_datos_6_bF_buf1_) );
BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[6]), .Y(bloque_datos_6_bF_buf0_) );
BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[68]), .Y(bloque_datos_68_bF_buf3_) );
BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[68]), .Y(bloque_datos_68_bF_buf2_) );
BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[68]), .Y(bloque_datos_68_bF_buf1_) );
BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[68]), .Y(bloque_datos_68_bF_buf0_) );
BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(_12844_), .Y(_12844__bF_buf4) );
BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(_12844_), .Y(_12844__bF_buf3) );
BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(_12844_), .Y(_12844__bF_buf2) );
BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(_12844_), .Y(_12844__bF_buf1) );
BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(_12844_), .Y(_12844__bF_buf0) );
BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[30]), .Y(bloque_datos_30_bF_buf3_) );
BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[30]), .Y(bloque_datos_30_bF_buf2_) );
BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[30]), .Y(bloque_datos_30_bF_buf1_) );
BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[30]), .Y(bloque_datos_30_bF_buf0_) );
BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[3]), .Y(bloque_datos_3_bF_buf3_) );
BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[3]), .Y(bloque_datos_3_bF_buf2_) );
BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[3]), .Y(bloque_datos_3_bF_buf1_) );
BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[3]), .Y(bloque_datos_3_bF_buf0_) );
BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[27]), .Y(bloque_datos_27_bF_buf4_) );
BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[27]), .Y(bloque_datos_27_bF_buf3_) );
BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[27]), .Y(bloque_datos_27_bF_buf2_) );
BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[27]), .Y(bloque_datos_27_bF_buf1_) );
BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[27]), .Y(bloque_datos_27_bF_buf0_) );
BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[65]), .Y(bloque_datos_65_bF_buf3_) );
BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[65]), .Y(bloque_datos_65_bF_buf2_) );
BUFX4 BUFX4_90 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[65]), .Y(bloque_datos_65_bF_buf1_) );
BUFX4 BUFX4_91 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[65]), .Y(bloque_datos_65_bF_buf0_) );
CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf10) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf9) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf8) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_9 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_10 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_11 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_92 ( .gnd(gnd), .vdd(vdd), .A(_4187_), .Y(_4187__bF_buf4) );
BUFX4 BUFX4_93 ( .gnd(gnd), .vdd(vdd), .A(_4187_), .Y(_4187__bF_buf3) );
BUFX4 BUFX4_94 ( .gnd(gnd), .vdd(vdd), .A(_4187_), .Y(_4187__bF_buf2) );
BUFX4 BUFX4_95 ( .gnd(gnd), .vdd(vdd), .A(_4187_), .Y(_4187__bF_buf1) );
BUFX4 BUFX4_96 ( .gnd(gnd), .vdd(vdd), .A(_4187_), .Y(_4187__bF_buf0) );
BUFX4 BUFX4_97 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[24]), .Y(bloque_datos_24_bF_buf4_) );
BUFX4 BUFX4_98 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[24]), .Y(bloque_datos_24_bF_buf3_) );
BUFX4 BUFX4_99 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[24]), .Y(bloque_datos_24_bF_buf2_) );
BUFX4 BUFX4_100 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[24]), .Y(bloque_datos_24_bF_buf1_) );
BUFX4 BUFX4_101 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[24]), .Y(bloque_datos_24_bF_buf0_) );
BUFX4 BUFX4_102 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[62]), .Y(bloque_datos_62_bF_buf3_) );
BUFX4 BUFX4_103 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[62]), .Y(bloque_datos_62_bF_buf2_) );
BUFX4 BUFX4_104 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[62]), .Y(bloque_datos_62_bF_buf1_) );
BUFX4 BUFX4_105 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[62]), .Y(bloque_datos_62_bF_buf0_) );
BUFX4 BUFX4_106 ( .gnd(gnd), .vdd(vdd), .A(_8323_), .Y(_8323__bF_buf3) );
BUFX4 BUFX4_107 ( .gnd(gnd), .vdd(vdd), .A(_8323_), .Y(_8323__bF_buf2) );
BUFX4 BUFX4_108 ( .gnd(gnd), .vdd(vdd), .A(_8323_), .Y(_8323__bF_buf1) );
BUFX4 BUFX4_109 ( .gnd(gnd), .vdd(vdd), .A(_8323_), .Y(_8323__bF_buf0) );
BUFX4 BUFX4_110 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[59]), .Y(bloque_datos_59_bF_buf4_) );
BUFX4 BUFX4_111 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[59]), .Y(bloque_datos_59_bF_buf3_) );
BUFX4 BUFX4_112 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[59]), .Y(bloque_datos_59_bF_buf2_) );
BUFX4 BUFX4_113 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[59]), .Y(bloque_datos_59_bF_buf1_) );
BUFX4 BUFX4_114 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[59]), .Y(bloque_datos_59_bF_buf0_) );
BUFX4 BUFX4_115 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[21]), .Y(bloque_datos_21_bF_buf3_) );
BUFX4 BUFX4_116 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[21]), .Y(bloque_datos_21_bF_buf2_) );
BUFX4 BUFX4_117 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[21]), .Y(bloque_datos_21_bF_buf1_) );
BUFX4 BUFX4_118 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[21]), .Y(bloque_datos_21_bF_buf0_) );
BUFX4 BUFX4_119 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[56]), .Y(bloque_datos_56_bF_buf4_) );
BUFX4 BUFX4_120 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[56]), .Y(bloque_datos_56_bF_buf3_) );
BUFX4 BUFX4_121 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[56]), .Y(bloque_datos_56_bF_buf2_) );
BUFX4 BUFX4_122 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[56]), .Y(bloque_datos_56_bF_buf1_) );
BUFX4 BUFX4_123 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[56]), .Y(bloque_datos_56_bF_buf0_) );
BUFX4 BUFX4_124 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[94]), .Y(bloque_datos_94_bF_buf3_) );
BUFX4 BUFX4_125 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[94]), .Y(bloque_datos_94_bF_buf2_) );
BUFX4 BUFX4_126 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[94]), .Y(bloque_datos_94_bF_buf1_) );
BUFX4 BUFX4_127 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[94]), .Y(bloque_datos_94_bF_buf0_) );
BUFX4 BUFX4_128 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[53]), .Y(bloque_datos_53_bF_buf3_) );
BUFX4 BUFX4_129 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[53]), .Y(bloque_datos_53_bF_buf2_) );
BUFX4 BUFX4_130 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[53]), .Y(bloque_datos_53_bF_buf1_) );
BUFX4 BUFX4_131 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[53]), .Y(bloque_datos_53_bF_buf0_) );
BUFX4 BUFX4_132 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[91]), .Y(bloque_datos_91_bF_buf3_) );
BUFX4 BUFX4_133 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[91]), .Y(bloque_datos_91_bF_buf2_) );
BUFX4 BUFX4_134 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[91]), .Y(bloque_datos_91_bF_buf1_) );
BUFX4 BUFX4_135 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[91]), .Y(bloque_datos_91_bF_buf0_) );
BUFX4 BUFX4_136 ( .gnd(gnd), .vdd(vdd), .A(_4234_), .Y(_4234__bF_buf4) );
BUFX4 BUFX4_137 ( .gnd(gnd), .vdd(vdd), .A(_4234_), .Y(_4234__bF_buf3) );
BUFX4 BUFX4_138 ( .gnd(gnd), .vdd(vdd), .A(_4234_), .Y(_4234__bF_buf2) );
BUFX4 BUFX4_139 ( .gnd(gnd), .vdd(vdd), .A(_4234_), .Y(_4234__bF_buf1) );
BUFX4 BUFX4_140 ( .gnd(gnd), .vdd(vdd), .A(_4234_), .Y(_4234__bF_buf0) );
BUFX4 BUFX4_141 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .Y(bloque_datos_88_bF_buf4_) );
BUFX4 BUFX4_142 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .Y(bloque_datos_88_bF_buf3_) );
BUFX4 BUFX4_143 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .Y(bloque_datos_88_bF_buf2_) );
BUFX4 BUFX4_144 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .Y(bloque_datos_88_bF_buf1_) );
BUFX4 BUFX4_145 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[88]), .Y(bloque_datos_88_bF_buf0_) );
BUFX4 BUFX4_146 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[12]), .Y(bloque_datos_12_bF_buf3_) );
BUFX4 BUFX4_147 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[12]), .Y(bloque_datos_12_bF_buf2_) );
BUFX4 BUFX4_148 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[12]), .Y(bloque_datos_12_bF_buf1_) );
BUFX4 BUFX4_149 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[12]), .Y(bloque_datos_12_bF_buf0_) );
BUFX4 BUFX4_150 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[50]), .Y(bloque_datos_50_bF_buf3_) );
BUFX4 BUFX4_151 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[50]), .Y(bloque_datos_50_bF_buf2_) );
BUFX4 BUFX4_152 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[50]), .Y(bloque_datos_50_bF_buf1_) );
BUFX4 BUFX4_153 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[50]), .Y(bloque_datos_50_bF_buf0_) );
BUFX4 BUFX4_154 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[47]), .Y(bloque_datos_47_bF_buf3_) );
BUFX4 BUFX4_155 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[47]), .Y(bloque_datos_47_bF_buf2_) );
BUFX4 BUFX4_156 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[47]), .Y(bloque_datos_47_bF_buf1_) );
BUFX4 BUFX4_157 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[47]), .Y(bloque_datos_47_bF_buf0_) );
BUFX4 BUFX4_158 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[85]), .Y(bloque_datos_85_bF_buf4_) );
BUFX4 BUFX4_159 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[85]), .Y(bloque_datos_85_bF_buf3_) );
BUFX4 BUFX4_160 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[85]), .Y(bloque_datos_85_bF_buf2_) );
BUFX4 BUFX4_161 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[85]), .Y(bloque_datos_85_bF_buf1_) );
BUFX4 BUFX4_162 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[85]), .Y(bloque_datos_85_bF_buf0_) );
BUFX4 BUFX4_163 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[44]), .Y(bloque_datos_44_bF_buf4_) );
BUFX4 BUFX4_164 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[44]), .Y(bloque_datos_44_bF_buf3_) );
BUFX4 BUFX4_165 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[44]), .Y(bloque_datos_44_bF_buf2_) );
BUFX4 BUFX4_166 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[44]), .Y(bloque_datos_44_bF_buf1_) );
BUFX4 BUFX4_167 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[44]), .Y(bloque_datos_44_bF_buf0_) );
BUFX4 BUFX4_168 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[82]), .Y(bloque_datos_82_bF_buf4_) );
BUFX4 BUFX4_169 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[82]), .Y(bloque_datos_82_bF_buf3_) );
BUFX4 BUFX4_170 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[82]), .Y(bloque_datos_82_bF_buf2_) );
BUFX4 BUFX4_171 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[82]), .Y(bloque_datos_82_bF_buf1_) );
BUFX4 BUFX4_172 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[82]), .Y(bloque_datos_82_bF_buf0_) );
BUFX4 BUFX4_173 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[79]), .Y(bloque_datos_79_bF_buf3_) );
BUFX4 BUFX4_174 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[79]), .Y(bloque_datos_79_bF_buf2_) );
BUFX4 BUFX4_175 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[79]), .Y(bloque_datos_79_bF_buf1_) );
BUFX4 BUFX4_176 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[79]), .Y(bloque_datos_79_bF_buf0_) );
BUFX4 BUFX4_177 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[41]), .Y(bloque_datos_41_bF_buf3_) );
BUFX4 BUFX4_178 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[41]), .Y(bloque_datos_41_bF_buf2_) );
BUFX4 BUFX4_179 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[41]), .Y(bloque_datos_41_bF_buf1_) );
BUFX4 BUFX4_180 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[41]), .Y(bloque_datos_41_bF_buf0_) );
BUFX4 BUFX4_181 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[38]), .Y(bloque_datos_38_bF_buf3_) );
BUFX4 BUFX4_182 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[38]), .Y(bloque_datos_38_bF_buf2_) );
BUFX4 BUFX4_183 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[38]), .Y(bloque_datos_38_bF_buf1_) );
BUFX4 BUFX4_184 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[38]), .Y(bloque_datos_38_bF_buf0_) );
BUFX4 BUFX4_185 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[76]), .Y(bloque_datos_76_bF_buf4_) );
BUFX4 BUFX4_186 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[76]), .Y(bloque_datos_76_bF_buf3_) );
BUFX4 BUFX4_187 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[76]), .Y(bloque_datos_76_bF_buf2_) );
BUFX4 BUFX4_188 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[76]), .Y(bloque_datos_76_bF_buf1_) );
BUFX4 BUFX4_189 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[76]), .Y(bloque_datos_76_bF_buf0_) );
BUFX4 BUFX4_190 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[35]), .Y(bloque_datos_35_bF_buf4_) );
BUFX4 BUFX4_191 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[35]), .Y(bloque_datos_35_bF_buf3_) );
BUFX4 BUFX4_192 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[35]), .Y(bloque_datos_35_bF_buf2_) );
BUFX4 BUFX4_193 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[35]), .Y(bloque_datos_35_bF_buf1_) );
BUFX4 BUFX4_194 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[35]), .Y(bloque_datos_35_bF_buf0_) );
BUFX4 BUFX4_195 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[73]), .Y(bloque_datos_73_bF_buf3_) );
BUFX4 BUFX4_196 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[73]), .Y(bloque_datos_73_bF_buf2_) );
BUFX4 BUFX4_197 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[73]), .Y(bloque_datos_73_bF_buf1_) );
BUFX4 BUFX4_198 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[73]), .Y(bloque_datos_73_bF_buf0_) );
BUFX4 BUFX4_199 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[32]), .Y(bloque_datos_32_bF_buf4_) );
BUFX4 BUFX4_200 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[32]), .Y(bloque_datos_32_bF_buf3_) );
BUFX4 BUFX4_201 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[32]), .Y(bloque_datos_32_bF_buf2_) );
BUFX4 BUFX4_202 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[32]), .Y(bloque_datos_32_bF_buf1_) );
BUFX4 BUFX4_203 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[32]), .Y(bloque_datos_32_bF_buf0_) );
BUFX4 BUFX4_204 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[70]), .Y(bloque_datos_70_bF_buf3_) );
BUFX4 BUFX4_205 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[70]), .Y(bloque_datos_70_bF_buf2_) );
BUFX4 BUFX4_206 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[70]), .Y(bloque_datos_70_bF_buf1_) );
BUFX4 BUFX4_207 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[70]), .Y(bloque_datos_70_bF_buf0_) );
BUFX4 BUFX4_208 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(inicio_bF_buf10) );
BUFX4 BUFX4_209 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(inicio_bF_buf9) );
BUFX4 BUFX4_210 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(inicio_bF_buf8) );
BUFX4 BUFX4_211 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(inicio_bF_buf7) );
BUFX4 BUFX4_212 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(inicio_bF_buf6) );
BUFX4 BUFX4_213 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(inicio_bF_buf5) );
BUFX4 BUFX4_214 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(inicio_bF_buf4) );
BUFX4 BUFX4_215 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(inicio_bF_buf3) );
BUFX4 BUFX4_216 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(inicio_bF_buf2) );
BUFX4 BUFX4_217 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(inicio_bF_buf1) );
BUFX4 BUFX4_218 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(inicio_bF_buf0) );
BUFX4 BUFX4_219 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[5]), .Y(bloque_datos_5_bF_buf3_) );
BUFX4 BUFX4_220 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[5]), .Y(bloque_datos_5_bF_buf2_) );
BUFX4 BUFX4_221 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[5]), .Y(bloque_datos_5_bF_buf1_) );
BUFX4 BUFX4_222 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[5]), .Y(bloque_datos_5_bF_buf0_) );
BUFX4 BUFX4_223 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[29]), .Y(bloque_datos_29_bF_buf4_) );
BUFX4 BUFX4_224 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[29]), .Y(bloque_datos_29_bF_buf3_) );
BUFX4 BUFX4_225 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[29]), .Y(bloque_datos_29_bF_buf2_) );
BUFX4 BUFX4_226 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[29]), .Y(bloque_datos_29_bF_buf1_) );
BUFX4 BUFX4_227 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[29]), .Y(bloque_datos_29_bF_buf0_) );
BUFX4 BUFX4_228 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[67]), .Y(bloque_datos_67_bF_buf4_) );
BUFX4 BUFX4_229 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[67]), .Y(bloque_datos_67_bF_buf3_) );
BUFX4 BUFX4_230 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[67]), .Y(bloque_datos_67_bF_buf2_) );
BUFX4 BUFX4_231 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[67]), .Y(bloque_datos_67_bF_buf1_) );
BUFX4 BUFX4_232 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[67]), .Y(bloque_datos_67_bF_buf0_) );
BUFX4 BUFX4_233 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[2]), .Y(bloque_datos_2_bF_buf3_) );
BUFX4 BUFX4_234 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[2]), .Y(bloque_datos_2_bF_buf2_) );
BUFX4 BUFX4_235 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[2]), .Y(bloque_datos_2_bF_buf1_) );
BUFX4 BUFX4_236 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[2]), .Y(bloque_datos_2_bF_buf0_) );
BUFX4 BUFX4_237 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[26]), .Y(bloque_datos_26_bF_buf3_) );
BUFX4 BUFX4_238 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[26]), .Y(bloque_datos_26_bF_buf2_) );
BUFX4 BUFX4_239 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[26]), .Y(bloque_datos_26_bF_buf1_) );
BUFX4 BUFX4_240 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[26]), .Y(bloque_datos_26_bF_buf0_) );
BUFX4 BUFX4_241 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[64]), .Y(bloque_datos_64_bF_buf4_) );
BUFX4 BUFX4_242 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[64]), .Y(bloque_datos_64_bF_buf3_) );
BUFX4 BUFX4_243 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[64]), .Y(bloque_datos_64_bF_buf2_) );
BUFX4 BUFX4_244 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[64]), .Y(bloque_datos_64_bF_buf1_) );
BUFX4 BUFX4_245 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[64]), .Y(bloque_datos_64_bF_buf0_) );
BUFX4 BUFX4_246 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[23]), .Y(bloque_datos_23_bF_buf3_) );
BUFX4 BUFX4_247 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[23]), .Y(bloque_datos_23_bF_buf2_) );
BUFX4 BUFX4_248 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[23]), .Y(bloque_datos_23_bF_buf1_) );
BUFX4 BUFX4_249 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[23]), .Y(bloque_datos_23_bF_buf0_) );
BUFX4 BUFX4_250 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[61]), .Y(bloque_datos_61_bF_buf4_) );
BUFX4 BUFX4_251 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[61]), .Y(bloque_datos_61_bF_buf3_) );
BUFX4 BUFX4_252 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[61]), .Y(bloque_datos_61_bF_buf2_) );
BUFX4 BUFX4_253 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[61]), .Y(bloque_datos_61_bF_buf1_) );
BUFX4 BUFX4_254 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[61]), .Y(bloque_datos_61_bF_buf0_) );
BUFX4 BUFX4_255 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[58]), .Y(bloque_datos_58_bF_buf4_) );
BUFX4 BUFX4_256 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[58]), .Y(bloque_datos_58_bF_buf3_) );
BUFX4 BUFX4_257 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[58]), .Y(bloque_datos_58_bF_buf2_) );
BUFX4 BUFX4_258 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[58]), .Y(bloque_datos_58_bF_buf1_) );
BUFX4 BUFX4_259 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[58]), .Y(bloque_datos_58_bF_buf0_) );
BUFX4 BUFX4_260 ( .gnd(gnd), .vdd(vdd), .A(_8492_), .Y(_8492__bF_buf4) );
BUFX4 BUFX4_261 ( .gnd(gnd), .vdd(vdd), .A(_8492_), .Y(_8492__bF_buf3) );
BUFX4 BUFX4_262 ( .gnd(gnd), .vdd(vdd), .A(_8492_), .Y(_8492__bF_buf2) );
BUFX4 BUFX4_263 ( .gnd(gnd), .vdd(vdd), .A(_8492_), .Y(_8492__bF_buf1) );
BUFX4 BUFX4_264 ( .gnd(gnd), .vdd(vdd), .A(_8492_), .Y(_8492__bF_buf0) );
BUFX4 BUFX4_265 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[20]), .Y(bloque_datos_20_bF_buf3_) );
BUFX4 BUFX4_266 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[20]), .Y(bloque_datos_20_bF_buf2_) );
BUFX4 BUFX4_267 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[20]), .Y(bloque_datos_20_bF_buf1_) );
BUFX4 BUFX4_268 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[20]), .Y(bloque_datos_20_bF_buf0_) );
BUFX4 BUFX4_269 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[93]), .Y(bloque_datos_93_bF_buf3_) );
BUFX4 BUFX4_270 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[93]), .Y(bloque_datos_93_bF_buf2_) );
BUFX4 BUFX4_271 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[93]), .Y(bloque_datos_93_bF_buf1_) );
BUFX4 BUFX4_272 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[93]), .Y(bloque_datos_93_bF_buf0_) );
BUFX4 BUFX4_273 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[14]), .Y(bloque_datos_14_bF_buf3_) );
BUFX4 BUFX4_274 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[14]), .Y(bloque_datos_14_bF_buf2_) );
BUFX4 BUFX4_275 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[14]), .Y(bloque_datos_14_bF_buf1_) );
BUFX4 BUFX4_276 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[14]), .Y(bloque_datos_14_bF_buf0_) );
BUFX4 BUFX4_277 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[52]), .Y(bloque_datos_52_bF_buf4_) );
BUFX4 BUFX4_278 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[52]), .Y(bloque_datos_52_bF_buf3_) );
BUFX4 BUFX4_279 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[52]), .Y(bloque_datos_52_bF_buf2_) );
BUFX4 BUFX4_280 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[52]), .Y(bloque_datos_52_bF_buf1_) );
BUFX4 BUFX4_281 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[52]), .Y(bloque_datos_52_bF_buf0_) );
BUFX4 BUFX4_282 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[90]), .Y(bloque_datos_90_bF_buf4_) );
BUFX4 BUFX4_283 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[90]), .Y(bloque_datos_90_bF_buf3_) );
BUFX4 BUFX4_284 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[90]), .Y(bloque_datos_90_bF_buf2_) );
BUFX4 BUFX4_285 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[90]), .Y(bloque_datos_90_bF_buf1_) );
BUFX4 BUFX4_286 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[90]), .Y(bloque_datos_90_bF_buf0_) );
BUFX4 BUFX4_287 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[49]), .Y(bloque_datos_49_bF_buf3_) );
BUFX4 BUFX4_288 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[49]), .Y(bloque_datos_49_bF_buf2_) );
BUFX4 BUFX4_289 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[49]), .Y(bloque_datos_49_bF_buf1_) );
BUFX4 BUFX4_290 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[49]), .Y(bloque_datos_49_bF_buf0_) );
BUFX4 BUFX4_291 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[87]), .Y(bloque_datos_87_bF_buf3_) );
BUFX4 BUFX4_292 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[87]), .Y(bloque_datos_87_bF_buf2_) );
BUFX4 BUFX4_293 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[87]), .Y(bloque_datos_87_bF_buf1_) );
BUFX4 BUFX4_294 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[87]), .Y(bloque_datos_87_bF_buf0_) );
BUFX4 BUFX4_295 ( .gnd(gnd), .vdd(vdd), .A(_8539_), .Y(_8539__bF_buf4) );
BUFX4 BUFX4_296 ( .gnd(gnd), .vdd(vdd), .A(_8539_), .Y(_8539__bF_buf3) );
BUFX4 BUFX4_297 ( .gnd(gnd), .vdd(vdd), .A(_8539_), .Y(_8539__bF_buf2) );
BUFX4 BUFX4_298 ( .gnd(gnd), .vdd(vdd), .A(_8539_), .Y(_8539__bF_buf1) );
BUFX4 BUFX4_299 ( .gnd(gnd), .vdd(vdd), .A(_8539_), .Y(_8539__bF_buf0) );
BUFX4 BUFX4_300 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[46]), .Y(bloque_datos_46_bF_buf4_) );
BUFX4 BUFX4_301 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[46]), .Y(bloque_datos_46_bF_buf3_) );
BUFX4 BUFX4_302 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[46]), .Y(bloque_datos_46_bF_buf2_) );
BUFX4 BUFX4_303 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[46]), .Y(bloque_datos_46_bF_buf1_) );
BUFX4 BUFX4_304 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[46]), .Y(bloque_datos_46_bF_buf0_) );
BUFX4 BUFX4_305 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[84]), .Y(bloque_datos_84_bF_buf4_) );
BUFX4 BUFX4_306 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[84]), .Y(bloque_datos_84_bF_buf3_) );
BUFX4 BUFX4_307 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[84]), .Y(bloque_datos_84_bF_buf2_) );
BUFX4 BUFX4_308 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[84]), .Y(bloque_datos_84_bF_buf1_) );
BUFX4 BUFX4_309 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[84]), .Y(bloque_datos_84_bF_buf0_) );
BUFX4 BUFX4_310 ( .gnd(gnd), .vdd(vdd), .A(_12628_), .Y(_12628__bF_buf3) );
BUFX4 BUFX4_311 ( .gnd(gnd), .vdd(vdd), .A(_12628_), .Y(_12628__bF_buf2) );
BUFX4 BUFX4_312 ( .gnd(gnd), .vdd(vdd), .A(_12628_), .Y(_12628__bF_buf1) );
BUFX4 BUFX4_313 ( .gnd(gnd), .vdd(vdd), .A(_12628_), .Y(_12628__bF_buf0) );
BUFX4 BUFX4_314 ( .gnd(gnd), .vdd(vdd), .A(_17149_), .Y(_17149__bF_buf4) );
BUFX4 BUFX4_315 ( .gnd(gnd), .vdd(vdd), .A(_17149_), .Y(_17149__bF_buf3) );
BUFX4 BUFX4_316 ( .gnd(gnd), .vdd(vdd), .A(_17149_), .Y(_17149__bF_buf2) );
BUFX4 BUFX4_317 ( .gnd(gnd), .vdd(vdd), .A(_17149_), .Y(_17149__bF_buf1) );
BUFX4 BUFX4_318 ( .gnd(gnd), .vdd(vdd), .A(_17149_), .Y(_17149__bF_buf0) );
BUFX4 BUFX4_319 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[43]), .Y(bloque_datos_43_bF_buf3_) );
BUFX4 BUFX4_320 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[43]), .Y(bloque_datos_43_bF_buf2_) );
BUFX4 BUFX4_321 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[43]), .Y(bloque_datos_43_bF_buf1_) );
BUFX4 BUFX4_322 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[43]), .Y(bloque_datos_43_bF_buf0_) );
BUFX4 BUFX4_323 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[81]), .Y(bloque_datos_81_bF_buf4_) );
BUFX4 BUFX4_324 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[81]), .Y(bloque_datos_81_bF_buf3_) );
BUFX4 BUFX4_325 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[81]), .Y(bloque_datos_81_bF_buf2_) );
BUFX4 BUFX4_326 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[81]), .Y(bloque_datos_81_bF_buf1_) );
BUFX4 BUFX4_327 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[81]), .Y(bloque_datos_81_bF_buf0_) );
BUFX4 BUFX4_328 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[78]), .Y(bloque_datos_78_bF_buf4_) );
BUFX4 BUFX4_329 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[78]), .Y(bloque_datos_78_bF_buf3_) );
BUFX4 BUFX4_330 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[78]), .Y(bloque_datos_78_bF_buf2_) );
BUFX4 BUFX4_331 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[78]), .Y(bloque_datos_78_bF_buf1_) );
BUFX4 BUFX4_332 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[78]), .Y(bloque_datos_78_bF_buf0_) );
BUFX4 BUFX4_333 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado), .Y(module_0_comparador_target_hash_0_terminado_bF_buf4) );
BUFX4 BUFX4_334 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado), .Y(module_0_comparador_target_hash_0_terminado_bF_buf3) );
BUFX4 BUFX4_335 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado), .Y(module_0_comparador_target_hash_0_terminado_bF_buf2) );
BUFX4 BUFX4_336 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado), .Y(module_0_comparador_target_hash_0_terminado_bF_buf1) );
BUFX4 BUFX4_337 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado), .Y(module_0_comparador_target_hash_0_terminado_bF_buf0) );
BUFX4 BUFX4_338 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[40]), .Y(bloque_datos_40_bF_buf4_) );
BUFX4 BUFX4_339 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[40]), .Y(bloque_datos_40_bF_buf3_) );
BUFX4 BUFX4_340 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[40]), .Y(bloque_datos_40_bF_buf2_) );
BUFX4 BUFX4_341 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[40]), .Y(bloque_datos_40_bF_buf1_) );
BUFX4 BUFX4_342 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[40]), .Y(bloque_datos_40_bF_buf0_) );
BUFX4 BUFX4_343 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado), .Y(module_2_comparador_target_hash_0_terminado_bF_buf6) );
BUFX4 BUFX4_344 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado), .Y(module_2_comparador_target_hash_0_terminado_bF_buf5) );
BUFX4 BUFX4_345 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado), .Y(module_2_comparador_target_hash_0_terminado_bF_buf4) );
BUFX4 BUFX4_346 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado), .Y(module_2_comparador_target_hash_0_terminado_bF_buf3) );
BUFX4 BUFX4_347 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado), .Y(module_2_comparador_target_hash_0_terminado_bF_buf2) );
BUFX4 BUFX4_348 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado), .Y(module_2_comparador_target_hash_0_terminado_bF_buf1) );
BUFX4 BUFX4_349 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado), .Y(module_2_comparador_target_hash_0_terminado_bF_buf0) );
BUFX4 BUFX4_350 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[37]), .Y(bloque_datos_37_bF_buf3_) );
BUFX4 BUFX4_351 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[37]), .Y(bloque_datos_37_bF_buf2_) );
BUFX4 BUFX4_352 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[37]), .Y(bloque_datos_37_bF_buf1_) );
BUFX4 BUFX4_353 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[37]), .Y(bloque_datos_37_bF_buf0_) );
BUFX4 BUFX4_354 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[75]), .Y(bloque_datos_75_bF_buf4_) );
BUFX4 BUFX4_355 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[75]), .Y(bloque_datos_75_bF_buf3_) );
BUFX4 BUFX4_356 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[75]), .Y(bloque_datos_75_bF_buf2_) );
BUFX4 BUFX4_357 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[75]), .Y(bloque_datos_75_bF_buf1_) );
BUFX4 BUFX4_358 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[75]), .Y(bloque_datos_75_bF_buf0_) );
BUFX4 BUFX4_359 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[34]), .Y(bloque_datos_34_bF_buf4_) );
BUFX4 BUFX4_360 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[34]), .Y(bloque_datos_34_bF_buf3_) );
BUFX4 BUFX4_361 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[34]), .Y(bloque_datos_34_bF_buf2_) );
BUFX4 BUFX4_362 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[34]), .Y(bloque_datos_34_bF_buf1_) );
BUFX4 BUFX4_363 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[34]), .Y(bloque_datos_34_bF_buf0_) );
BUFX4 BUFX4_364 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[72]), .Y(bloque_datos_72_bF_buf4_) );
BUFX4 BUFX4_365 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[72]), .Y(bloque_datos_72_bF_buf3_) );
BUFX4 BUFX4_366 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[72]), .Y(bloque_datos_72_bF_buf2_) );
BUFX4 BUFX4_367 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[72]), .Y(bloque_datos_72_bF_buf1_) );
BUFX4 BUFX4_368 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[72]), .Y(bloque_datos_72_bF_buf0_) );
BUFX4 BUFX4_369 ( .gnd(gnd), .vdd(vdd), .A(_17102_), .Y(_17102__bF_buf4) );
BUFX4 BUFX4_370 ( .gnd(gnd), .vdd(vdd), .A(_17102_), .Y(_17102__bF_buf3) );
BUFX4 BUFX4_371 ( .gnd(gnd), .vdd(vdd), .A(_17102_), .Y(_17102__bF_buf2) );
BUFX4 BUFX4_372 ( .gnd(gnd), .vdd(vdd), .A(_17102_), .Y(_17102__bF_buf1) );
BUFX4 BUFX4_373 ( .gnd(gnd), .vdd(vdd), .A(_17102_), .Y(_17102__bF_buf0) );
BUFX4 BUFX4_374 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[69]), .Y(bloque_datos_69_bF_buf3_) );
BUFX4 BUFX4_375 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[69]), .Y(bloque_datos_69_bF_buf2_) );
BUFX4 BUFX4_376 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[69]), .Y(bloque_datos_69_bF_buf1_) );
BUFX4 BUFX4_377 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[69]), .Y(bloque_datos_69_bF_buf0_) );
BUFX4 BUFX4_378 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[31]), .Y(bloque_datos_31_bF_buf3_) );
BUFX4 BUFX4_379 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[31]), .Y(bloque_datos_31_bF_buf2_) );
BUFX4 BUFX4_380 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[31]), .Y(bloque_datos_31_bF_buf1_) );
BUFX4 BUFX4_381 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[31]), .Y(bloque_datos_31_bF_buf0_) );
BUFX4 BUFX4_382 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[4]), .Y(bloque_datos_4_bF_buf3_) );
BUFX4 BUFX4_383 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[4]), .Y(bloque_datos_4_bF_buf2_) );
BUFX4 BUFX4_384 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[4]), .Y(bloque_datos_4_bF_buf1_) );
BUFX4 BUFX4_385 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[4]), .Y(bloque_datos_4_bF_buf0_) );
BUFX4 BUFX4_386 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[28]), .Y(bloque_datos_28_bF_buf4_) );
BUFX4 BUFX4_387 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[28]), .Y(bloque_datos_28_bF_buf3_) );
BUFX4 BUFX4_388 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[28]), .Y(bloque_datos_28_bF_buf2_) );
BUFX4 BUFX4_389 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[28]), .Y(bloque_datos_28_bF_buf1_) );
BUFX4 BUFX4_390 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[28]), .Y(bloque_datos_28_bF_buf0_) );
BUFX4 BUFX4_391 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[66]), .Y(bloque_datos_66_bF_buf4_) );
BUFX4 BUFX4_392 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[66]), .Y(bloque_datos_66_bF_buf3_) );
BUFX4 BUFX4_393 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[66]), .Y(bloque_datos_66_bF_buf2_) );
BUFX4 BUFX4_394 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[66]), .Y(bloque_datos_66_bF_buf1_) );
BUFX4 BUFX4_395 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[66]), .Y(bloque_datos_66_bF_buf0_) );
BUFX4 BUFX4_396 ( .gnd(gnd), .vdd(vdd), .A(_4018_), .Y(_4018__bF_buf3) );
BUFX4 BUFX4_397 ( .gnd(gnd), .vdd(vdd), .A(_4018_), .Y(_4018__bF_buf2) );
BUFX4 BUFX4_398 ( .gnd(gnd), .vdd(vdd), .A(_4018_), .Y(_4018__bF_buf1) );
BUFX4 BUFX4_399 ( .gnd(gnd), .vdd(vdd), .A(_4018_), .Y(_4018__bF_buf0) );
BUFX4 BUFX4_400 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[25]), .Y(bloque_datos_25_bF_buf3_) );
BUFX4 BUFX4_401 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[25]), .Y(bloque_datos_25_bF_buf2_) );
BUFX4 BUFX4_402 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[25]), .Y(bloque_datos_25_bF_buf1_) );
BUFX4 BUFX4_403 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[25]), .Y(bloque_datos_25_bF_buf0_) );
BUFX4 BUFX4_404 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[22]), .Y(bloque_datos_22_bF_buf3_) );
BUFX4 BUFX4_405 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[22]), .Y(bloque_datos_22_bF_buf2_) );
BUFX4 BUFX4_406 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[22]), .Y(bloque_datos_22_bF_buf1_) );
BUFX4 BUFX4_407 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[22]), .Y(bloque_datos_22_bF_buf0_) );
BUFX4 BUFX4_408 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[60]), .Y(bloque_datos_60_bF_buf3_) );
BUFX4 BUFX4_409 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[60]), .Y(bloque_datos_60_bF_buf2_) );
BUFX4 BUFX4_410 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[60]), .Y(bloque_datos_60_bF_buf1_) );
BUFX4 BUFX4_411 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[60]), .Y(bloque_datos_60_bF_buf0_) );
BUFX4 BUFX4_412 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[19]), .Y(bloque_datos_19_bF_buf3_) );
BUFX4 BUFX4_413 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[19]), .Y(bloque_datos_19_bF_buf2_) );
BUFX4 BUFX4_414 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[19]), .Y(bloque_datos_19_bF_buf1_) );
BUFX4 BUFX4_415 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[19]), .Y(bloque_datos_19_bF_buf0_) );
BUFX4 BUFX4_416 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[57]), .Y(bloque_datos_57_bF_buf3_) );
BUFX4 BUFX4_417 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[57]), .Y(bloque_datos_57_bF_buf2_) );
BUFX4 BUFX4_418 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[57]), .Y(bloque_datos_57_bF_buf1_) );
BUFX4 BUFX4_419 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[57]), .Y(bloque_datos_57_bF_buf0_) );
BUFX4 BUFX4_420 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[95]), .Y(bloque_datos_95_bF_buf3_) );
BUFX4 BUFX4_421 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[95]), .Y(bloque_datos_95_bF_buf2_) );
BUFX4 BUFX4_422 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[95]), .Y(bloque_datos_95_bF_buf1_) );
BUFX4 BUFX4_423 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[95]), .Y(bloque_datos_95_bF_buf0_) );
BUFX4 BUFX4_424 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[16]), .Y(bloque_datos_16_bF_buf3_) );
BUFX4 BUFX4_425 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[16]), .Y(bloque_datos_16_bF_buf2_) );
BUFX4 BUFX4_426 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[16]), .Y(bloque_datos_16_bF_buf1_) );
BUFX4 BUFX4_427 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[16]), .Y(bloque_datos_16_bF_buf0_) );
BUFX4 BUFX4_428 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[54]), .Y(bloque_datos_54_bF_buf3_) );
BUFX4 BUFX4_429 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[54]), .Y(bloque_datos_54_bF_buf2_) );
BUFX4 BUFX4_430 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[54]), .Y(bloque_datos_54_bF_buf1_) );
BUFX4 BUFX4_431 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[54]), .Y(bloque_datos_54_bF_buf0_) );
BUFX4 BUFX4_432 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[92]), .Y(bloque_datos_92_bF_buf3_) );
BUFX4 BUFX4_433 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[92]), .Y(bloque_datos_92_bF_buf2_) );
BUFX4 BUFX4_434 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[92]), .Y(bloque_datos_92_bF_buf1_) );
BUFX4 BUFX4_435 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[92]), .Y(bloque_datos_92_bF_buf0_) );
BUFX4 BUFX4_436 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[89]), .Y(bloque_datos_89_bF_buf3_) );
BUFX4 BUFX4_437 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[89]), .Y(bloque_datos_89_bF_buf2_) );
BUFX4 BUFX4_438 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[89]), .Y(bloque_datos_89_bF_buf1_) );
BUFX4 BUFX4_439 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[89]), .Y(bloque_datos_89_bF_buf0_) );
BUFX4 BUFX4_440 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[13]), .Y(bloque_datos_13_bF_buf3_) );
BUFX4 BUFX4_441 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[13]), .Y(bloque_datos_13_bF_buf2_) );
BUFX4 BUFX4_442 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[13]), .Y(bloque_datos_13_bF_buf1_) );
BUFX4 BUFX4_443 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[13]), .Y(bloque_datos_13_bF_buf0_) );
BUFX4 BUFX4_444 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[51]), .Y(bloque_datos_51_bF_buf4_) );
BUFX4 BUFX4_445 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[51]), .Y(bloque_datos_51_bF_buf3_) );
BUFX4 BUFX4_446 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[51]), .Y(bloque_datos_51_bF_buf2_) );
BUFX4 BUFX4_447 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[51]), .Y(bloque_datos_51_bF_buf1_) );
BUFX4 BUFX4_448 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[51]), .Y(bloque_datos_51_bF_buf0_) );
BUFX4 BUFX4_449 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[48]), .Y(bloque_datos_48_bF_buf4_) );
BUFX4 BUFX4_450 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[48]), .Y(bloque_datos_48_bF_buf3_) );
BUFX4 BUFX4_451 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[48]), .Y(bloque_datos_48_bF_buf2_) );
BUFX4 BUFX4_452 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[48]), .Y(bloque_datos_48_bF_buf1_) );
BUFX4 BUFX4_453 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[48]), .Y(bloque_datos_48_bF_buf0_) );
BUFX4 BUFX4_454 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[86]), .Y(bloque_datos_86_bF_buf4_) );
BUFX4 BUFX4_455 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[86]), .Y(bloque_datos_86_bF_buf3_) );
BUFX4 BUFX4_456 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[86]), .Y(bloque_datos_86_bF_buf2_) );
BUFX4 BUFX4_457 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[86]), .Y(bloque_datos_86_bF_buf1_) );
BUFX4 BUFX4_458 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[86]), .Y(bloque_datos_86_bF_buf0_) );
BUFX4 BUFX4_459 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[45]), .Y(bloque_datos_45_bF_buf4_) );
BUFX4 BUFX4_460 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[45]), .Y(bloque_datos_45_bF_buf3_) );
BUFX4 BUFX4_461 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[45]), .Y(bloque_datos_45_bF_buf2_) );
BUFX4 BUFX4_462 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[45]), .Y(bloque_datos_45_bF_buf1_) );
BUFX4 BUFX4_463 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[45]), .Y(bloque_datos_45_bF_buf0_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_0__0_), .Y(bounty_out[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_0__1_), .Y(bounty_out[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_0__2_), .Y(bounty_out[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_0__3_), .Y(bounty_out[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(bounty_out[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(bounty_out[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(bounty_out[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(bounty_out[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(bounty_out[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(bounty_out[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(bounty_out[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(bounty_out[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(bounty_out[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(bounty_out[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(bounty_out[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(bounty_out[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(bounty_out[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(bounty_out[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(bounty_out[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(bounty_out[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(bounty_out[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(bounty_out[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(bounty_out[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(bounty_out[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(terminado_out) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(bounty_72_), .B(module_3_comparador_target_hash_0_terminado_bF_buf1), .Y(_2_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf2), .B(bounty_0_), .Y(_3_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(bounty_24_), .B(module_1_comparador_target_hash_0_terminado_bF_buf5), .C(module_2_comparador_target_hash_0_terminado_bF_buf6), .Y(_4_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(module_1_comparador_target_hash_0_terminado_bF_buf5), .C(_4_), .Y(_5_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(bounty_48_), .Y(_6_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf4), .B(_6_), .C(module_3_comparador_target_hash_0_terminado_bF_buf0), .Y(_7_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_5_), .Y(_8_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(_8_), .Y(_0__0_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf1), .B(bounty_73_), .Y(_9_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf0), .B(bounty_1_), .Y(_10_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf6), .B(bounty_25_), .C(module_2_comparador_target_hash_0_terminado_bF_buf5), .Y(_11_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(module_1_comparador_target_hash_0_terminado_bF_buf6), .C(_11_), .Y(_12_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(bounty_49_), .Y(_13_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf4), .B(_13_), .C(module_3_comparador_target_hash_0_terminado_bF_buf0), .Y(_14_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_12_), .Y(_15_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_15_), .Y(_0__1_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf1), .B(bounty_74_), .Y(_16_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_2_), .Y(_17_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_26_), .C(module_2_comparador_target_hash_0_terminado_bF_buf1), .Y(_18_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(module_1_comparador_target_hash_0_terminado_bF_buf4), .C(_18_), .Y(_19_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(bounty_50_), .Y(_20_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf4), .B(_20_), .C(module_3_comparador_target_hash_0_terminado_bF_buf0), .Y(_21_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_19_), .Y(_22_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_22_), .Y(_0__2_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf1), .B(bounty_75_), .Y(_23_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_3_), .Y(_24_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf5), .B(bounty_27_), .C(module_2_comparador_target_hash_0_terminado_bF_buf6), .Y(_25_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(module_1_comparador_target_hash_0_terminado_bF_buf0), .C(_25_), .Y(_26_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(bounty_51_), .Y(_27_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf2), .B(_27_), .C(module_3_comparador_target_hash_0_terminado_bF_buf0), .Y(_28_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_26_), .Y(_29_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_29_), .Y(_0__3_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf1), .B(bounty_76_), .Y(_30_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_4_), .Y(_31_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf6), .B(bounty_28_), .C(module_2_comparador_target_hash_0_terminado_bF_buf5), .Y(_32_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(module_1_comparador_target_hash_0_terminado_bF_buf1), .C(_32_), .Y(_33_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(bounty_52_), .Y(_34_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf4), .B(_34_), .C(module_3_comparador_target_hash_0_terminado_bF_buf0), .Y(_35_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_33_), .Y(_36_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_36_), .Y(_0__4_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf1), .B(bounty_77_), .Y(_37_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf0), .B(bounty_5_), .Y(_38_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf6), .B(bounty_29_), .C(module_2_comparador_target_hash_0_terminado_bF_buf5), .Y(_39_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(module_1_comparador_target_hash_0_terminado_bF_buf1), .C(_39_), .Y(_40_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(bounty_53_), .Y(_41_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf2), .B(_41_), .C(module_3_comparador_target_hash_0_terminado_bF_buf2), .Y(_42_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_40_), .Y(_43_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_43_), .Y(_0__5_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_78_), .Y(_44_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf0), .B(bounty_6_), .Y(_45_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf0), .B(bounty_30_), .C(module_2_comparador_target_hash_0_terminado_bF_buf5), .Y(_46_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(module_1_comparador_target_hash_0_terminado_bF_buf1), .C(_46_), .Y(_47_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(bounty_54_), .Y(_48_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf2), .B(_48_), .C(module_3_comparador_target_hash_0_terminado_bF_buf2), .Y(_49_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_47_), .Y(_50_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_50_), .Y(_0__6_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_79_), .Y(_51_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf2), .B(bounty_7_), .Y(_52_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf5), .B(bounty_31_), .C(module_2_comparador_target_hash_0_terminado_bF_buf6), .Y(_53_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(module_1_comparador_target_hash_0_terminado_bF_buf5), .C(_53_), .Y(_54_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(bounty_55_), .Y(_55_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf2), .B(_55_), .C(module_3_comparador_target_hash_0_terminado_bF_buf2), .Y(_56_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_54_), .Y(_57_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_57_), .Y(_0__7_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_80_), .Y(_58_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf1), .B(bounty_8_), .Y(_59_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf2), .B(bounty_32_), .C(module_2_comparador_target_hash_0_terminado_bF_buf0), .Y(_60_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(module_1_comparador_target_hash_0_terminado_bF_buf2), .C(_60_), .Y(_61_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(bounty_56_), .Y(_62_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf0), .B(_62_), .C(module_3_comparador_target_hash_0_terminado_bF_buf4), .Y(_63_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_61_), .Y(_64_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_64_), .Y(_0__8_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_81_), .Y(_65_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_9_), .Y(_66_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf2), .B(bounty_33_), .C(module_2_comparador_target_hash_0_terminado_bF_buf0), .Y(_67_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(module_1_comparador_target_hash_0_terminado_bF_buf2), .C(_67_), .Y(_68_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(bounty_57_), .Y(_69_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf3), .B(_69_), .C(module_3_comparador_target_hash_0_terminado_bF_buf5), .Y(_70_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_68_), .Y(_71_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_71_), .Y(_0__9_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf6), .B(bounty_82_), .Y(_72_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf1), .B(bounty_10_), .Y(_73_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_34_), .C(module_2_comparador_target_hash_0_terminado_bF_buf1), .Y(_74_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(module_1_comparador_target_hash_0_terminado_bF_buf3), .C(_74_), .Y(_75_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(bounty_58_), .Y(_76_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf3), .B(_76_), .C(module_3_comparador_target_hash_0_terminado_bF_buf6), .Y(_77_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_75_), .Y(_78_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_78_), .Y(_0__10_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_83_), .Y(_79_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf1), .B(bounty_11_), .Y(_80_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf2), .B(bounty_35_), .C(module_2_comparador_target_hash_0_terminado_bF_buf0), .Y(_81_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(module_1_comparador_target_hash_0_terminado_bF_buf2), .C(_81_), .Y(_82_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(bounty_59_), .Y(_83_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf0), .B(_83_), .C(module_3_comparador_target_hash_0_terminado_bF_buf6), .Y(_84_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_82_), .Y(_85_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_85_), .Y(_0__11_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_84_), .Y(_86_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_12_), .Y(_87_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf5), .B(bounty_36_), .C(module_2_comparador_target_hash_0_terminado_bF_buf6), .Y(_88_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(module_1_comparador_target_hash_0_terminado_bF_buf0), .C(_88_), .Y(_89_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(bounty_60_), .Y(_90_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf2), .B(_90_), .C(module_3_comparador_target_hash_0_terminado_bF_buf5), .Y(_91_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_89_), .Y(_92_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_92_), .Y(_0__12_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf2), .B(bounty_85_), .Y(_93_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_13_), .Y(_94_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf1), .B(bounty_37_), .C(module_2_comparador_target_hash_0_terminado_bF_buf5), .Y(_95_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(module_1_comparador_target_hash_0_terminado_bF_buf1), .C(_95_), .Y(_96_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(bounty_61_), .Y(_97_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf2), .B(_97_), .C(module_3_comparador_target_hash_0_terminado_bF_buf2), .Y(_98_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_96_), .Y(_99_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_99_), .Y(_0__13_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf2), .B(bounty_86_), .Y(_100_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_14_), .Y(_101_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf5), .B(bounty_38_), .C(module_2_comparador_target_hash_0_terminado_bF_buf6), .Y(_102_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(module_1_comparador_target_hash_0_terminado_bF_buf1), .C(_102_), .Y(_103_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(bounty_62_), .Y(_104_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf4), .B(_104_), .C(module_3_comparador_target_hash_0_terminado_bF_buf0), .Y(_105_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_103_), .Y(_106_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_106_), .Y(_0__14_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf1), .B(bounty_87_), .Y(_107_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf2), .B(bounty_15_), .Y(_108_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf0), .B(bounty_39_), .C(module_2_comparador_target_hash_0_terminado_bF_buf6), .Y(_109_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(module_1_comparador_target_hash_0_terminado_bF_buf0), .C(_109_), .Y(_110_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(bounty_63_), .Y(_111_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf4), .B(_111_), .C(module_3_comparador_target_hash_0_terminado_bF_buf0), .Y(_112_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_110_), .Y(_113_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_113_), .Y(_0__15_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_88_), .Y(_114_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_16_), .Y(_115_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_40_), .C(module_2_comparador_target_hash_0_terminado_bF_buf1), .Y(_116_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(module_1_comparador_target_hash_0_terminado_bF_buf4), .C(_116_), .Y(_117_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(bounty_64_), .Y(_118_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf0), .B(_118_), .C(module_3_comparador_target_hash_0_terminado_bF_buf6), .Y(_119_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_117_), .Y(_120_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_120_), .Y(_0__16_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_89_), .Y(_121_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_17_), .Y(_122_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_41_), .C(module_2_comparador_target_hash_0_terminado_bF_buf1), .Y(_123_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(module_1_comparador_target_hash_0_terminado_bF_buf3), .C(_123_), .Y(_124_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(bounty_65_), .Y(_125_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf3), .B(_125_), .C(module_3_comparador_target_hash_0_terminado_bF_buf6), .Y(_126_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_124_), .Y(_127_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_127_), .Y(_0__17_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_90_), .Y(_128_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_18_), .Y(_129_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_42_), .C(module_2_comparador_target_hash_0_terminado_bF_buf1), .Y(_130_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(module_1_comparador_target_hash_0_terminado_bF_buf3), .C(_130_), .Y(_131_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(bounty_66_), .Y(_132_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf3), .B(_132_), .C(module_3_comparador_target_hash_0_terminado_bF_buf5), .Y(_133_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_131_), .Y(_134_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_134_), .Y(_0__18_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_91_), .Y(_135_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf1), .B(bounty_19_), .Y(_136_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_43_), .C(module_2_comparador_target_hash_0_terminado_bF_buf1), .Y(_137_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(module_1_comparador_target_hash_0_terminado_bF_buf3), .C(_137_), .Y(_138_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(bounty_67_), .Y(_139_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf3), .B(_139_), .C(module_3_comparador_target_hash_0_terminado_bF_buf6), .Y(_140_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_138_), .Y(_141_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_141_), .Y(_0__19_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_92_), .Y(_142_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf2), .B(bounty_20_), .Y(_143_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_44_), .C(module_2_comparador_target_hash_0_terminado_bF_buf1), .Y(_144_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(module_1_comparador_target_hash_0_terminado_bF_buf4), .C(_144_), .Y(_145_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(bounty_68_), .Y(_146_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf2), .B(_146_), .C(module_3_comparador_target_hash_0_terminado_bF_buf5), .Y(_147_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_145_), .Y(_148_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_148_), .Y(_0__20_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf2), .B(bounty_93_), .Y(_149_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf2), .B(bounty_21_), .Y(_150_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf6), .B(bounty_45_), .C(module_2_comparador_target_hash_0_terminado_bF_buf5), .Y(_151_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(module_1_comparador_target_hash_0_terminado_bF_buf6), .C(_151_), .Y(_152_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(bounty_69_), .Y(_153_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf3), .B(_153_), .C(module_3_comparador_target_hash_0_terminado_bF_buf5), .Y(_154_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_152_), .Y(_155_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_155_), .Y(_0__21_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf3), .B(bounty_94_), .Y(_156_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf0), .B(bounty_22_), .Y(_157_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf0), .B(bounty_46_), .C(module_2_comparador_target_hash_0_terminado_bF_buf6), .Y(_158_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(module_1_comparador_target_hash_0_terminado_bF_buf0), .C(_158_), .Y(_159_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(bounty_70_), .Y(_160_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf4), .B(_160_), .C(module_3_comparador_target_hash_0_terminado_bF_buf5), .Y(_161_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_159_), .Y(_162_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_162_), .Y(_0__22_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(module_3_comparador_target_hash_0_terminado_bF_buf4), .B(bounty_95_), .Y(_163_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf0), .B(bounty_23_), .Y(_164_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(module_1_comparador_target_hash_0_terminado_bF_buf6), .B(bounty_47_), .C(module_2_comparador_target_hash_0_terminado_bF_buf5), .Y(_165_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(module_1_comparador_target_hash_0_terminado_bF_buf1), .C(_165_), .Y(_166_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(bounty_71_), .Y(_167_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf3), .B(_167_), .C(module_3_comparador_target_hash_0_terminado_bF_buf5), .Y(_168_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_166_), .Y(_169_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_169_), .Y(_0__23_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(module_0_comparador_target_hash_0_terminado_bF_buf1), .B(module_1_comparador_target_hash_0_terminado_bF_buf2), .Y(_170_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(module_2_comparador_target_hash_0_terminado_bF_buf0), .B(module_3_comparador_target_hash_0_terminado_bF_buf6), .Y(_171_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_171_), .Y(_1_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_405_), .C(_406_), .Y(_407_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_200_), .B(_389_), .Y(_408_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(module_0_W_200_), .Y(_409_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_409_), .Y(_410_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_410_), .C(_402_), .Y(_411_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_402_), .Y(_412_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(_410_), .Y(_413_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_412_), .C(_2395_), .Y(_414_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_228_), .B(_411_), .C(_414_), .Y(_415_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_228_), .Y(_416_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_406_), .C(_404_), .Y(_417_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_3824_), .B(_397_), .C(_394_), .Y(_418_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_3827_), .B(_399_), .C(_400_), .Y(_419_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_419_), .C(_3880_), .Y(_420_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_420_), .C(_413_), .Y(_421_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_2384_), .B(_411_), .C(_421_), .Y(_422_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_422_), .Y(_423_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_415_), .C(_3836_), .Y(_424_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_3836_), .Y(_425_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_228_), .B(_422_), .Y(_426_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_411_), .C(_414_), .Y(_427_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_427_), .C(_425_), .Y(_428_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_428_), .C(_3878_), .Y(_429_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_3842_), .B(_3844_), .C(_3837_), .Y(_430_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_426_), .C(_427_), .Y(_431_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3836_), .B(_423_), .C(_415_), .Y(_432_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_431_), .C(_432_), .Y(_433_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_216_), .B(_410_), .Y(_434_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(module_0_W_216_), .Y(_435_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_435_), .Y(_436_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_436_), .C(_429_), .Y(_437_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_432_), .C(_430_), .Y(_438_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_428_), .C(_3878_), .Y(_439_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(_436_), .Y(_440_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_438_), .C(_440_), .Y(_441_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_3629_), .B(_437_), .C(_441_), .Y(_442_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_244_), .B(_442_), .Y(_443_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_244_), .Y(_444_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_429_), .Y(_445_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_445_), .C(_3630_), .Y(_446_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_437_), .C(_446_), .Y(_447_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_3877_), .B(_447_), .C(_443_), .Y(_448_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_244_), .B(_437_), .C(_446_), .Y(_449_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_442_), .Y(_450_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_3849_), .B(_449_), .C(_450_), .Y(_451_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_448_), .B(_451_), .C(_3876_), .Y(_452_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_3625_), .B(_3850_), .Y(_453_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_3640_), .B(_3853_), .C(_453_), .Y(_454_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_450_), .C(_3849_), .Y(_455_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_443_), .C(_3877_), .Y(_456_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_454_), .C(_456_), .Y(_457_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_232_), .B(_440_), .Y(_458_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(module_0_W_232_), .Y(_459_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_459_), .Y(_460_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_452_), .C(_460_), .Y(_461_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_456_), .C(_454_), .Y(_462_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_448_), .B(_451_), .C(_3876_), .Y(_463_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(_460_), .Y(_464_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_463_), .C(_462_), .Y(_465_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_461_), .Y(_466_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_3873_), .Y(module_0_H_4_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_3873_), .B(_465_), .C(_461_), .Y(_467_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_216_), .B(_413_), .Y(_468_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_200_), .B(_390_), .Y(_469_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_184_), .B(_365_), .Y(_470_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_343_), .Y(_471_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_168_), .B(_471_), .Y(_472_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_152_), .B(_321_), .Y(_473_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_153_), .Y(_474_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_136_), .B(_298_), .Y(_475_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_137_), .Y(_476_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_268_), .Y(_477_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf4_), .B(_477_), .Y(_478_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf3_), .Y(_479_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_73_bF_buf3_), .Y(_480_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf4_), .B(_218_), .Y(_481_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf4_), .B(_193_), .Y(_482_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf4_), .B(_3979_), .Y(_483_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .B(_3954_), .Y(_484_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_25_), .Y(_485_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_9_), .Y(_486_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_486_), .Y(_487_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_25_), .B(module_0_W_9_), .Y(_488_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_487_), .Y(_489_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_3952_), .B(_489_), .Y(_490_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_3952_), .Y(_491_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_491_), .Y(_492_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .B(_492_), .Y(_493_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .Y(_494_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_490_), .Y(_495_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_495_), .Y(_496_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_493_), .C(_484_), .Y(_497_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_493_), .Y(_498_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_484_), .Y(_499_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_497_), .Y(_500_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf3_), .B(_500_), .Y(_501_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(bloque_datos_25_bF_buf2_), .Y(_502_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_501_), .C(_483_), .Y(_503_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_501_), .Y(_504_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_504_), .B(_483_), .Y(_505_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_503_), .Y(_506_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf3_), .B(_506_), .Y(_507_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf2_), .Y(_508_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_505_), .Y(_509_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_509_), .Y(_510_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_510_), .C(_482_), .Y(_511_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_510_), .Y(_512_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_482_), .Y(_513_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_511_), .Y(_514_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf3_), .B(_514_), .Y(_515_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf2_), .Y(_516_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_511_), .B(_513_), .Y(_517_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_517_), .Y(_518_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_518_), .C(_481_), .Y(_519_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_518_), .Y(_520_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_481_), .Y(_521_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_521_), .Y(_522_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_522_), .Y(_523_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_480_), .Y(_524_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_524_), .Y(_525_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_525_), .Y(_526_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(_265_), .Y(_527_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_527_), .Y(_528_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_528_), .Y(_529_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_479_), .Y(_530_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_530_), .Y(_531_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_531_), .Y(_532_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_531_), .Y(_533_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_533_), .Y(_534_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_532_), .B(_534_), .Y(_535_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_535_), .Y(_536_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(_535_), .Y(_537_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_137_), .B(_537_), .Y(_538_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_538_), .Y(_539_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_539_), .Y(_540_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_539_), .Y(_541_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_541_), .Y(_542_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_542_), .Y(_543_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_543_), .Y(_544_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_543_), .Y(_545_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_545_), .Y(_546_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_546_), .Y(_547_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_547_), .Y(_548_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_547_), .Y(_549_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_549_), .Y(_550_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_550_), .Y(_551_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(_551_), .Y(_552_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_169_), .B(_552_), .Y(_553_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_169_), .B(_552_), .Y(_554_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(_554_), .Y(_555_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_555_), .B(_553_), .C(_472_), .Y(_556_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(_555_), .Y(_557_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_168_), .B(_471_), .C(_557_), .Y(_558_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_558_), .Y(_559_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(_559_), .Y(_560_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_185_), .B(_560_), .Y(_561_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_185_), .B(_560_), .Y(_562_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(_562_), .Y(_563_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_561_), .C(_470_), .Y(_564_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_563_), .Y(_565_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_184_), .B(_365_), .C(_565_), .Y(_566_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_564_), .B(_566_), .Y(_567_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(_567_), .Y(_568_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_201_), .B(_568_), .Y(_569_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_201_), .B(_568_), .Y(_570_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(_570_), .Y(_571_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_569_), .C(_469_), .Y(_572_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_571_), .Y(_573_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_200_), .B(_390_), .C(_573_), .Y(_574_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_574_), .Y(_575_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(_575_), .Y(_576_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_217_), .B(_576_), .Y(_577_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_217_), .B(_576_), .Y(_578_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(_578_), .Y(_579_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_577_), .C(_468_), .Y(_580_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_579_), .Y(_581_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_216_), .B(_413_), .C(_581_), .Y(_582_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_582_), .Y(_583_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(_583_), .Y(_584_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_233_), .B(_584_), .Y(_585_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_233_), .B(_584_), .Y(_586_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(_586_), .Y(_587_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_585_), .C(_458_), .Y(_588_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_587_), .Y(_589_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_232_), .B(_440_), .C(_589_), .Y(_590_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_590_), .Y(_591_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_454_), .C(_448_), .Y(_592_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_245_), .Y(_593_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_432_), .C(_424_), .Y(_594_) );
INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(_426_), .Y(_595_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_229_), .Y(_596_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_406_), .C(_398_), .Y(_597_) );
INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(_399_), .Y(_598_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_213_), .Y(_599_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_382_), .C(_374_), .Y(_600_) );
INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(_378_), .Y(_601_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_197_), .Y(_602_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_356_), .C(_351_), .Y(_603_) );
INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(_352_), .Y(_604_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_181_), .Y(_605_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_3886_), .B(_339_), .C(_332_), .Y(_606_) );
INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(_334_), .Y(_607_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_165_), .Y(_608_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_543_), .Y(_609_) );
AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_314_), .C(_307_), .Y(_610_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_308_), .Y(_611_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_149_), .Y(_612_) );
AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_3889_), .C(_294_), .Y(_613_) );
AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_258_), .C(_3891_), .Y(_614_) );
AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_263_), .C(_614_), .Y(_615_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_3743_), .C(_229_), .Y(_616_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_616_), .B(_3893_), .C(_238_), .Y(_617_) );
AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_208_), .C(_3897_), .Y(_618_) );
AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_211_), .C(_618_), .Y(_619_) );
AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_183_), .C(_3901_), .Y(_620_) );
AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_186_), .C(_620_), .Y(_621_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_3972_), .Y(_622_) );
AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_3971_), .B(_3973_), .C(_622_), .Y(_623_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_3948_), .Y(_624_) );
AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_3949_), .B(_3947_), .C(_624_), .Y(_625_) );
AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_3921_), .B(_3920_), .C(_3680_), .Y(_626_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_3932_), .Y(_627_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_3920_), .Y(_628_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_2779_), .B(_2768_), .Y(_629_) );
INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_5_), .Y(_630_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_3912_), .B(_630_), .Y(_631_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_631_), .Y(_632_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_629_), .Y(_633_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_5_), .B(_3912_), .Y(_634_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_630_), .B(_3909_), .Y(_635_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_634_), .C(_633_), .Y(_636_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_21_), .B(_632_), .C(_636_), .Y(_637_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_21_), .Y(_638_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_634_), .C(_629_), .Y(_639_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .B(_2779_), .C(_631_), .Y(_640_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_640_), .C(_639_), .Y(_641_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_637_), .C(_641_), .Y(_642_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_21_), .B(_640_), .C(_639_), .Y(_643_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_632_), .C(_636_), .Y(_644_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_3920_), .B(_644_), .C(_643_), .Y(_645_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_645_), .Y(_646_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_646_), .B(_627_), .Y(_647_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_642_), .Y(_648_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_3932_), .C(_648_), .Y(_649_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_2855_), .B(module_0_W_9_), .Y(_650_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_649_), .C(_647_), .Y(_651_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_3919_), .B(_3923_), .Y(_652_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_652_), .Y(_653_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_646_), .B(_627_), .Y(_654_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_650_), .Y(_655_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_653_), .C(_655_), .Y(_656_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf3_), .B(_651_), .C(_656_), .Y(_657_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf2_), .Y(_658_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_649_), .C(_647_), .Y(_659_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_653_), .C(_650_), .Y(_660_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_659_), .C(_660_), .Y(_661_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_657_), .C(_661_), .Y(_662_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf1_), .B(_659_), .C(_660_), .Y(_663_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_651_), .C(_656_), .Y(_664_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_3941_), .B(_663_), .C(_664_), .Y(_665_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_625_), .B(_662_), .C(_665_), .Y(_666_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_3948_), .B(_3950_), .Y(_667_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_3941_), .B(_657_), .C(_661_), .Y(_668_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_663_), .C(_664_), .Y(_669_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_669_), .C(_667_), .Y(_670_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_2899_), .B(_492_), .Y(_671_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_671_), .Y(_672_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_672_), .C(_670_), .Y(_673_) );
AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_669_), .C(_667_), .Y(_674_) );
AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_665_), .C(_625_), .Y(_675_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_675_), .C(_671_), .Y(_676_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf3_), .B(_673_), .C(_676_), .Y(_677_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf2_), .Y(_678_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_671_), .C(_670_), .Y(_679_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_675_), .C(_672_), .Y(_680_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_679_), .C(_680_), .Y(_681_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_3961_), .B(_677_), .C(_681_), .Y(_682_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf1_), .B(_679_), .C(_680_), .Y(_683_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_673_), .C(_676_), .Y(_684_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_3967_), .B(_683_), .C(_684_), .Y(_685_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_682_), .B(_685_), .C(_623_), .Y(_686_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_3973_), .Y(_687_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(_3902_), .C(_3972_), .Y(_688_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_3967_), .B(_677_), .C(_681_), .Y(_689_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_3961_), .B(_683_), .C(_684_), .Y(_690_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_688_), .C(_690_), .Y(_691_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_499_), .Y(_692_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_2954_), .B(_692_), .Y(_693_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_693_), .Y(_694_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_691_), .C(_686_), .Y(_695_) );
AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_690_), .C(_688_), .Y(_696_) );
AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_682_), .B(_685_), .C(_623_), .Y(_697_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_697_), .C(_693_), .Y(_698_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf3_), .B(_695_), .C(_698_), .Y(_699_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf2_), .Y(_700_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_691_), .C(_686_), .Y(_701_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_697_), .C(_694_), .Y(_702_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_701_), .C(_702_), .Y(_703_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_699_), .C(_703_), .Y(_704_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf1_), .B(_701_), .C(_702_), .Y(_705_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_695_), .C(_698_), .Y(_706_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_705_), .C(_706_), .Y(_707_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_704_), .C(_707_), .Y(_708_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_3719_), .C(_180_), .Y(_709_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_3900_), .C(_187_), .Y(_710_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_699_), .C(_703_), .Y(_711_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_705_), .C(_706_), .Y(_712_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_710_), .B(_711_), .C(_712_), .Y(_713_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_3031_), .B(_506_), .Y(_714_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_708_), .C(_713_), .Y(_715_) );
AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_712_), .C(_710_), .Y(_716_) );
AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_707_), .C(_621_), .Y(_717_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_714_), .Y(_718_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_717_), .C(_718_), .Y(_719_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf3_), .B(_715_), .C(_719_), .Y(_720_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf2_), .Y(_721_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_708_), .C(_713_), .Y(_722_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_717_), .C(_714_), .Y(_723_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_721_), .B(_722_), .C(_723_), .Y(_724_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_720_), .C(_724_), .Y(_725_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf1_), .B(_722_), .C(_723_), .Y(_726_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_721_), .B(_715_), .C(_719_), .Y(_727_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_726_), .C(_727_), .Y(_728_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_725_), .C(_728_), .Y(_729_) );
NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_206_), .C(_204_), .Y(_730_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_730_), .B(_3895_), .C(_212_), .Y(_731_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_720_), .C(_724_), .Y(_732_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_726_), .C(_727_), .Y(_733_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_733_), .C(_731_), .Y(_734_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3097_), .B(_514_), .Y(_735_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_735_), .Y(_736_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_736_), .B(_729_), .C(_734_), .Y(_737_) );
AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_733_), .C(_731_), .Y(_738_) );
AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(_728_), .C(_619_), .Y(_739_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_738_), .B(_739_), .C(_735_), .Y(_740_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf3_), .B(_737_), .C(_740_), .Y(_741_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf2_), .Y(_742_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_729_), .C(_734_), .Y(_743_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_738_), .B(_739_), .C(_736_), .Y(_744_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_742_), .B(_743_), .C(_744_), .Y(_745_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_741_), .C(_745_), .Y(_746_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf1_), .B(_743_), .C(_744_), .Y(_747_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_742_), .B(_737_), .C(_740_), .Y(_748_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_747_), .C(_748_), .Y(_749_) );
AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_749_), .C(_617_), .Y(_750_) );
AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_232_), .C(_3894_), .Y(_751_) );
AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_239_), .C(_751_), .Y(_752_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_741_), .C(_745_), .Y(_753_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_747_), .C(_748_), .Y(_754_) );
AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_754_), .C(_752_), .Y(_755_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_3141_), .B(_522_), .Y(_756_) );
NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_756_), .C(_750_), .Y(_757_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_753_), .C(_754_), .Y(_758_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_749_), .C(_617_), .Y(_759_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_756_), .Y(_760_) );
AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(_759_), .C(_760_), .Y(_761_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_757_), .B(_761_), .C(bloque_datos_85_bF_buf4_), .Y(_762_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf3_), .Y(_763_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_760_), .B(_758_), .C(_759_), .Y(_764_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_755_), .C(_756_), .Y(_765_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_763_), .B(_764_), .C(_765_), .Y(_766_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_766_), .C(_762_), .Y(_767_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf2_), .B(_764_), .C(_765_), .Y(_768_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_757_), .B(_761_), .C(_763_), .Y(_769_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_768_), .C(_769_), .Y(_770_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_767_), .C(_770_), .Y(_771_) );
NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_3755_), .C(_255_), .Y(_772_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_3890_), .C(_262_), .Y(_773_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_766_), .C(_762_), .Y(_774_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_768_), .C(_769_), .Y(_775_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_774_), .B(_775_), .C(_773_), .Y(_776_) );
XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3239_), .B(_528_), .Y(_777_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_771_), .C(_776_), .Y(_778_) );
AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_774_), .B(_775_), .C(_773_), .Y(_779_) );
AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_770_), .C(_615_), .Y(_780_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_777_), .Y(_781_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_779_), .B(_780_), .C(_781_), .Y(_782_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_133_), .B(_778_), .C(_782_), .Y(_783_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_133_), .Y(_784_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_781_), .B(_771_), .C(_776_), .Y(_785_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_779_), .B(_780_), .C(_777_), .Y(_786_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_784_), .B(_785_), .C(_786_), .Y(_787_) );
AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_787_), .C(_275_), .Y(_788_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_133_), .B(_785_), .C(_786_), .Y(_789_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_784_), .B(_778_), .C(_782_), .Y(_790_) );
AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_790_), .C(_282_), .Y(_791_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_791_), .C(_613_), .Y(_792_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_286_), .C(_280_), .Y(_793_) );
AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_787_), .C(_282_), .Y(_794_) );
AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_790_), .C(_275_), .Y(_795_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_795_), .C(_793_), .Y(_796_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_792_), .C(_796_), .Y(_797_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_789_), .C(_790_), .Y(_798_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_783_), .C(_787_), .Y(_799_) );
AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_799_), .C(_793_), .Y(_800_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_789_), .C(_790_), .Y(_801_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_783_), .C(_787_), .Y(_802_) );
AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_801_), .B(_802_), .C(_613_), .Y(_803_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_803_), .C(_535_), .Y(_804_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(_804_), .Y(_805_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_612_), .B(_3316_), .C(_805_), .Y(_806_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_803_), .C(_537_), .Y(_807_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_792_), .C(_796_), .Y(_808_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_3316_), .B(_808_), .C(_807_), .Y(_809_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_149_), .B(_809_), .Y(_810_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_806_), .C(_810_), .Y(_811_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_149_), .B(_809_), .Y(_812_) );
AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_3316_), .B(_805_), .C(_612_), .Y(_813_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_813_), .C(_308_), .Y(_814_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_811_), .B(_610_), .C(_814_), .Y(_815_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_3888_), .C(_313_), .Y(_816_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_813_), .C(_611_), .Y(_817_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_806_), .C(_810_), .Y(_818_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_817_), .C(_816_), .Y(_819_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_815_), .C(_819_), .Y(_820_) );
AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_817_), .C(_816_), .Y(_821_) );
AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_811_), .B(_814_), .C(_610_), .Y(_822_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_821_), .B(_822_), .C(_543_), .Y(_823_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_820_), .B(_823_), .Y(_824_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(_3400_), .C(_824_), .Y(_825_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_821_), .B(_822_), .C(_609_), .Y(_826_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_815_), .C(_819_), .Y(_827_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_3400_), .B(_827_), .C(_826_), .Y(_828_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_165_), .B(_828_), .Y(_829_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_825_), .C(_829_), .Y(_830_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_165_), .B(_828_), .Y(_831_) );
AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_3400_), .B(_824_), .C(_608_), .Y(_832_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_831_), .B(_832_), .C(_334_), .Y(_833_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_830_), .C(_833_), .Y(_834_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_3887_), .B(_336_), .C(_338_), .Y(_835_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_831_), .B(_832_), .C(_607_), .Y(_836_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_825_), .C(_829_), .Y(_837_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_837_), .B(_835_), .C(_836_), .Y(_838_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_834_), .C(_838_), .Y(_839_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_834_), .B(_838_), .Y(_840_) );
AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_840_), .C(_3409_), .Y(_841_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_839_), .C(_841_), .Y(_842_) );
AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_837_), .B(_836_), .C(_835_), .Y(_843_) );
AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_830_), .B(_833_), .C(_606_), .Y(_844_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_844_), .C(_552_), .Y(_845_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .B(_839_), .C(_845_), .Y(_846_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_181_), .B(_846_), .Y(_847_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_842_), .C(_847_), .Y(_848_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_181_), .B(_846_), .Y(_849_) );
AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_841_), .C(_605_), .Y(_850_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_849_), .B(_850_), .C(_352_), .Y(_851_) );
NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_848_), .C(_851_), .Y(_852_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_3884_), .C(_357_), .Y(_853_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_849_), .B(_850_), .C(_604_), .Y(_854_) );
NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_842_), .C(_847_), .Y(_855_) );
NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_853_), .C(_854_), .Y(_856_) );
NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(_852_), .C(_856_), .Y(_857_) );
AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_854_), .C(_853_), .Y(_858_) );
AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_851_), .C(_603_), .Y(_859_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_858_), .B(_859_), .C(_559_), .Y(_860_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_857_), .B(_860_), .Y(_861_) );
NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(_3417_), .C(_861_), .Y(_862_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_858_), .B(_859_), .C(_560_), .Y(_863_) );
NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_852_), .C(_856_), .Y(_864_) );
NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_3417_), .B(_864_), .C(_863_), .Y(_865_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_197_), .B(_865_), .Y(_866_) );
NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(_862_), .C(_866_), .Y(_867_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_197_), .B(_865_), .Y(_868_) );
AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_3417_), .B(_861_), .C(_602_), .Y(_869_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_869_), .C(_378_), .Y(_870_) );
NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_600_), .C(_870_), .Y(_871_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_3882_), .C(_383_), .Y(_872_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_869_), .C(_601_), .Y(_873_) );
NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_862_), .C(_866_), .Y(_874_) );
NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(_874_), .B(_873_), .C(_872_), .Y(_875_) );
NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_871_), .C(_875_), .Y(_876_) );
AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_874_), .B(_873_), .C(_872_), .Y(_877_) );
AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_870_), .C(_600_), .Y(_878_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_877_), .B(_878_), .C(_567_), .Y(_879_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_876_), .B(_879_), .Y(_880_) );
NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_599_), .B(_3425_), .C(_880_), .Y(_881_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_877_), .B(_878_), .C(_568_), .Y(_882_) );
NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_871_), .C(_875_), .Y(_883_) );
NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_3425_), .B(_883_), .C(_882_), .Y(_884_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_213_), .B(_884_), .Y(_885_) );
NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_881_), .C(_885_), .Y(_886_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_213_), .B(_884_), .Y(_887_) );
AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_3425_), .B(_880_), .C(_599_), .Y(_888_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_887_), .B(_888_), .C(_399_), .Y(_889_) );
NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_597_), .C(_889_), .Y(_890_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_3880_), .C(_405_), .Y(_891_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_887_), .B(_888_), .C(_598_), .Y(_892_) );
NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_881_), .C(_885_), .Y(_893_) );
NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_891_), .C(_892_), .Y(_894_) );
NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_576_), .B(_890_), .C(_894_), .Y(_895_) );
AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_892_), .C(_891_), .Y(_896_) );
AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_889_), .C(_597_), .Y(_897_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_896_), .B(_897_), .C(_575_), .Y(_898_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_895_), .B(_898_), .Y(_899_) );
NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_3434_), .C(_899_), .Y(_900_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_896_), .B(_897_), .C(_576_), .Y(_901_) );
NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_890_), .C(_894_), .Y(_902_) );
NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_3434_), .B(_902_), .C(_901_), .Y(_903_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_229_), .B(_903_), .Y(_904_) );
NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_900_), .C(_904_), .Y(_905_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_229_), .B(_903_), .Y(_906_) );
AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_3434_), .B(_899_), .C(_596_), .Y(_907_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_906_), .B(_907_), .C(_426_), .Y(_908_) );
NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_905_), .C(_908_), .Y(_909_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_3878_), .B(_428_), .C(_431_), .Y(_910_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_906_), .B(_907_), .C(_595_), .Y(_911_) );
NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_900_), .C(_904_), .Y(_912_) );
NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_912_), .C(_911_), .Y(_913_) );
NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_909_), .C(_913_), .Y(_914_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_913_), .Y(_915_) );
AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_915_), .C(_3631_), .Y(_916_) );
NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_914_), .C(_916_), .Y(_917_) );
AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_912_), .B(_911_), .C(_910_), .Y(_918_) );
AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_908_), .C(_594_), .Y(_919_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_918_), .B(_919_), .C(_584_), .Y(_920_) );
NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_3442_), .B(_914_), .C(_920_), .Y(_921_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_245_), .B(_921_), .Y(_922_) );
NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_917_), .C(_922_), .Y(_923_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_443_), .Y(_924_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_245_), .B(_921_), .Y(_925_) );
AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_914_), .B(_916_), .C(_593_), .Y(_926_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_925_), .B(_926_), .C(_924_), .Y(_927_) );
NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_592_), .C(_927_), .Y(_928_) );
AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_3876_), .C(_455_), .Y(_929_) );
NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_924_), .B(_926_), .C(_925_), .Y(_930_) );
AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_922_), .C(_443_), .Y(_931_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_931_), .C(_929_), .Y(_932_) );
NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_928_), .C(_932_), .Y(_933_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_591_), .Y(_934_) );
NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_929_), .C(_927_), .Y(_935_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_931_), .C(_592_), .Y(_936_) );
NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_935_), .C(_936_), .Y(_937_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_937_), .Y(_938_) );
XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_467_), .Y(module_0_H_5_) );
AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_937_), .C(_467_), .Y(_939_) );
AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_592_), .C(_931_), .Y(_940_) );
AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_900_), .B(_904_), .C(_426_), .Y(_941_) );
AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_912_), .B(_910_), .C(_941_), .Y(_942_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_3612_), .Y(_943_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_3613_), .Y(_944_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(_943_), .Y(_945_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_945_), .Y(_946_) );
AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_885_), .C(_399_), .Y(_947_) );
AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_891_), .C(_947_), .Y(_948_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_3602_), .Y(_949_) );
AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_866_), .C(_378_), .Y(_950_) );
AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_874_), .B(_872_), .C(_950_), .Y(_951_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_3592_), .B(_3591_), .Y(_952_) );
INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(_952_), .Y(_953_) );
NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_850_), .C(_849_), .Y(_954_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_954_), .B(_603_), .C(_854_), .Y(_955_) );
INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(_3584_), .Y(_956_) );
AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_829_), .C(_334_), .Y(_957_) );
AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_837_), .B(_835_), .C(_957_), .Y(_958_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_817_), .Y(_959_) );
AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_816_), .C(_959_), .Y(_960_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_3563_), .B(_3564_), .Y(_961_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_961_), .Y(_962_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_791_), .B(_613_), .C(_798_), .Y(_963_) );
INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(_789_), .Y(_964_) );
AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_762_), .C(_257_), .Y(_965_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_965_), .B(_615_), .C(_774_), .Y(_966_) );
INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(_762_), .Y(_967_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_759_), .Y(_968_) );
INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(_741_), .Y(_969_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_734_), .Y(_970_) );
INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(_720_), .Y(_971_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_713_), .Y(_972_) );
INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(_699_), .Y(_973_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_691_), .Y(_974_) );
INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(_677_), .Y(_975_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_669_), .Y(_976_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_625_), .C(_668_), .Y(_977_) );
INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(_657_), .Y(_978_) );
NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_3920_), .B(_637_), .C(_641_), .Y(_979_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_637_), .Y(_980_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_3459_), .B(_3463_), .Y(_981_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_981_), .Y(_982_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_6_), .Y(_983_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_983_), .Y(_984_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_634_), .Y(_985_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_984_), .B(_985_), .C(_982_), .Y(_986_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_985_), .B(_984_), .Y(_987_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_3460_), .B(_3461_), .C(_987_), .Y(_988_) );
NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_22_), .B(_986_), .C(_988_), .Y(_989_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_22_), .Y(_990_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_984_), .B(_985_), .C(_981_), .Y(_991_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_987_), .Y(_992_) );
NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_991_), .C(_992_), .Y(_993_) );
NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(_980_), .B(_993_), .C(_989_), .Y(_994_) );
AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_991_), .B(_992_), .C(_990_), .Y(_995_) );
AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_986_), .B(_988_), .C(module_0_W_22_), .Y(_996_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_995_), .C(_637_), .Y(_997_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_997_), .Y(_998_) );
AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_979_), .B(_649_), .C(_998_), .Y(_999_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_999_), .Y(_1000_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_646_), .C(_979_), .Y(_1001_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_998_), .Y(_1002_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_1002_), .B(_1001_), .Y(_1003_) );
INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_10_), .Y(_1004_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .B(_3470_), .Y(_1005_) );
XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .B(_1004_), .Y(_1006_) );
NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .B(_1006_), .C(_1003_), .Y(_1007_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .B(_1002_), .Y(_1008_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .Y(_1009_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_999_), .C(_1009_), .Y(_1010_) );
NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf3_), .B(_1010_), .C(_1007_), .Y(_1011_) );
INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf2_), .Y(_1012_) );
NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .B(_1009_), .C(_1003_), .Y(_1013_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_999_), .C(_1006_), .Y(_1014_) );
NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1012_), .B(_1014_), .C(_1013_), .Y(_1015_) );
NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_1011_), .C(_1015_), .Y(_1016_) );
NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf1_), .B(_1014_), .C(_1013_), .Y(_1017_) );
NAND3X1 NAND3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1012_), .B(_1010_), .C(_1007_), .Y(_1018_) );
NAND3X1 NAND3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_1017_), .C(_1018_), .Y(_1019_) );
NAND3X1 NAND3X1_172 ( .gnd(gnd), .vdd(vdd), .A(_977_), .B(_1016_), .C(_1019_), .Y(_1020_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_668_), .Y(_1021_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1021_), .B(_675_), .Y(_1022_) );
AOI21X1 AOI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .B(_1018_), .C(_657_), .Y(_1023_) );
AOI21X1 AOI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(_1015_), .C(_978_), .Y(_1024_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(_1024_), .C(_1022_), .Y(_1025_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_3482_), .B(_3489_), .Y(_1026_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_26_), .B(module_0_W_10_), .Y(_1027_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_26_), .Y(_1028_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_1004_), .Y(_1029_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(_1027_), .Y(_1030_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_1030_), .Y(_1031_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .B(_1029_), .Y(_1032_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_486_), .C(_1032_), .Y(_1033_) );
NAND3X1 NAND3X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .B(_1033_), .C(_491_), .Y(_1034_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_24_), .B(module_0_W_8_), .C(_489_), .Y(_1035_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_487_), .Y(_1036_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1036_), .B(_1032_), .Y(_1037_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_1030_), .Y(_1038_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1038_), .B(_1037_), .C(_1035_), .Y(_1039_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1034_), .Y(_1040_) );
XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .B(_1040_), .Y(_1041_) );
NAND3X1 NAND3X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_1041_), .C(_1025_), .Y(_1042_) );
NAND3X1 NAND3X1_175 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_1011_), .C(_1015_), .Y(_1043_) );
NAND3X1 NAND3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_1017_), .C(_1018_), .Y(_1044_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_670_), .C(_1043_), .D(_1044_), .Y(_1045_) );
AOI21X1 AOI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_1019_), .C(_977_), .Y(_1046_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .Y(_1047_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(_1046_), .C(_1047_), .Y(_1048_) );
NAND3X1 NAND3X1_177 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf3_), .B(_1042_), .C(_1048_), .Y(_1049_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf2_), .Y(_1050_) );
NAND3X1 NAND3X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_1047_), .C(_1025_), .Y(_1051_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(_1046_), .C(_1041_), .Y(_1052_) );
NAND3X1 NAND3X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1050_), .B(_1051_), .C(_1052_), .Y(_1053_) );
NAND3X1 NAND3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_975_), .B(_1049_), .C(_1053_), .Y(_1054_) );
NAND3X1 NAND3X1_181 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf1_), .B(_1051_), .C(_1052_), .Y(_1055_) );
NAND3X1 NAND3X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1050_), .B(_1042_), .C(_1048_), .Y(_1056_) );
NAND3X1 NAND3X1_183 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_1055_), .C(_1056_), .Y(_1057_) );
NAND3X1 NAND3X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1054_), .B(_1057_), .C(_974_), .Y(_1058_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_691_), .B(_689_), .Y(_1059_) );
AOI21X1 AOI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1056_), .C(_677_), .Y(_1060_) );
AOI21X1 AOI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_1053_), .C(_975_), .Y(_1061_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1060_), .B(_1061_), .C(_1059_), .Y(_1062_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_3499_), .B(_3496_), .Y(_1063_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(_498_), .Y(_1064_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_496_), .Y(_1065_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .Y(_1066_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_1040_), .Y(_1067_) );
NAND3X1 NAND3X1_185 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .B(_1039_), .C(_1034_), .Y(_1068_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1067_), .Y(_1069_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1065_), .B(_1069_), .Y(_1070_) );
AOI21X1 AOI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1067_), .C(_496_), .Y(_1071_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1071_), .B(_1070_), .Y(_1072_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1064_), .B(_1072_), .Y(_1073_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .B(_1071_), .C(_499_), .Y(_1074_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1074_), .B(_1073_), .Y(_1075_) );
XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .B(_1075_), .Y(_1076_) );
NAND3X1 NAND3X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .B(_1076_), .C(_1062_), .Y(_1077_) );
NAND3X1 NAND3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_1049_), .C(_1053_), .Y(_1078_) );
NAND3X1 NAND3X1_188 ( .gnd(gnd), .vdd(vdd), .A(_975_), .B(_1055_), .C(_1056_), .Y(_1079_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_691_), .C(_1078_), .D(_1079_), .Y(_1080_) );
AOI21X1 AOI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1054_), .B(_1057_), .C(_974_), .Y(_1081_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_1076_), .Y(_1082_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1081_), .C(_1082_), .Y(_1083_) );
NAND3X1 NAND3X1_189 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf3_), .B(_1083_), .C(_1077_), .Y(_1084_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf2_), .Y(_1085_) );
NAND3X1 NAND3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .B(_1082_), .C(_1062_), .Y(_1086_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1081_), .C(_1076_), .Y(_1087_) );
NAND3X1 NAND3X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1085_), .B(_1087_), .C(_1086_), .Y(_1088_) );
NAND3X1 NAND3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_973_), .B(_1084_), .C(_1088_), .Y(_1089_) );
NAND3X1 NAND3X1_193 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf1_), .B(_1087_), .C(_1086_), .Y(_1090_) );
NAND3X1 NAND3X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1085_), .B(_1083_), .C(_1077_), .Y(_1091_) );
NAND3X1 NAND3X1_195 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_1090_), .C(_1091_), .Y(_1092_) );
NAND3X1 NAND3X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_1092_), .C(_972_), .Y(_1093_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_711_), .Y(_1094_) );
AOI21X1 AOI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1091_), .C(_699_), .Y(_1095_) );
AOI21X1 AOI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_1088_), .C(_973_), .Y(_1096_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_1096_), .C(_1094_), .Y(_1097_) );
INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf3_), .Y(_1098_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_1064_), .Y(_1099_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_1074_), .Y(_1100_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1099_), .B(_1100_), .C(_1098_), .Y(_1101_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_1075_), .B(_1098_), .Y(_1102_) );
NAND3X1 NAND3X1_197 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_1101_), .C(_1102_), .Y(_1103_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_502_), .Y(_1104_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .Y(_1105_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1098_), .B(_1075_), .Y(_1106_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(_1106_), .C(_1104_), .Y(_1107_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1103_), .B(_1107_), .Y(_1108_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_1108_), .B(_505_), .Y(_1109_) );
NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .B(_1106_), .C(_1105_), .Y(_1110_) );
AOI21X1 AOI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .B(_1102_), .C(_502_), .Y(_1111_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1110_), .B(_1111_), .C(_505_), .Y(_1112_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1112_), .B(_1109_), .Y(_1113_) );
XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_3728_), .B(_1113_), .Y(_1114_) );
NAND3X1 NAND3X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .B(_1114_), .C(_1097_), .Y(_1115_) );
NAND3X1 NAND3X1_199 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_1084_), .C(_1088_), .Y(_1116_) );
NAND3X1 NAND3X1_200 ( .gnd(gnd), .vdd(vdd), .A(_973_), .B(_1090_), .C(_1091_), .Y(_1117_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_713_), .C(_1116_), .D(_1117_), .Y(_1118_) );
AOI21X1 AOI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_1092_), .C(_972_), .Y(_1119_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(_1114_), .Y(_1120_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1118_), .B(_1119_), .C(_1120_), .Y(_1121_) );
NAND3X1 NAND3X1_201 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf3_), .B(_1115_), .C(_1121_), .Y(_1122_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf2_), .Y(_1123_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1118_), .B(_1119_), .C(_1114_), .Y(_1124_) );
NAND3X1 NAND3X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .B(_1120_), .C(_1097_), .Y(_1125_) );
NAND3X1 NAND3X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_1125_), .C(_1124_), .Y(_1126_) );
NAND3X1 NAND3X1_204 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_1122_), .C(_1126_), .Y(_1127_) );
NAND3X1 NAND3X1_205 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf1_), .B(_1125_), .C(_1124_), .Y(_1128_) );
NAND3X1 NAND3X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_1115_), .C(_1121_), .Y(_1129_) );
NAND3X1 NAND3X1_207 ( .gnd(gnd), .vdd(vdd), .A(_720_), .B(_1128_), .C(_1129_), .Y(_1130_) );
NAND3X1 NAND3X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .B(_1130_), .C(_970_), .Y(_1131_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_732_), .Y(_1132_) );
AOI21X1 AOI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(_1129_), .C(_720_), .Y(_1133_) );
AOI21X1 AOI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .B(_1126_), .C(_971_), .Y(_1134_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .B(_1134_), .C(_1132_), .Y(_1135_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(_510_), .Y(_1136_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf3_), .Y(_1137_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_1108_), .Y(_1138_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_1112_), .Y(_1139_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1139_), .B(_1138_), .C(_1137_), .Y(_1140_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .Y(_1141_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_1113_), .Y(_1142_) );
NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_1136_), .C(_1142_), .Y(_1143_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(_1139_), .Y(_1144_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf2_), .B(_1144_), .Y(_1145_) );
AOI21X1 AOI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1145_), .C(_510_), .Y(_1146_) );
NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_1146_), .C(_1143_), .Y(_1147_) );
INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(_513_), .Y(_1148_) );
NAND3X1 NAND3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_1140_), .C(_1145_), .Y(_1149_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .B(_1141_), .C(_1136_), .Y(_1150_) );
AOI21X1 AOI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1149_), .B(_1150_), .C(_1148_), .Y(_1151_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1151_), .B(_1147_), .Y(_1152_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_3519_), .B(_3520_), .C(_1152_), .Y(_1153_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_3520_), .B(_3519_), .Y(_1154_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1151_), .C(_1154_), .Y(_1155_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1155_), .Y(_1156_) );
NAND3X1 NAND3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1131_), .B(_1156_), .C(_1135_), .Y(_1157_) );
NAND3X1 NAND3X1_211 ( .gnd(gnd), .vdd(vdd), .A(_720_), .B(_1122_), .C(_1126_), .Y(_1158_) );
NAND3X1 NAND3X1_212 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_1128_), .C(_1129_), .Y(_1159_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_734_), .C(_1158_), .D(_1159_), .Y(_1160_) );
AOI21X1 AOI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .B(_1130_), .C(_970_), .Y(_1161_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_1156_), .Y(_1162_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_1161_), .C(_1162_), .Y(_1163_) );
NAND3X1 NAND3X1_213 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf3_), .B(_1157_), .C(_1163_), .Y(_1164_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf2_), .Y(_1165_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_1161_), .C(_1156_), .Y(_1166_) );
NAND3X1 NAND3X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1131_), .B(_1162_), .C(_1135_), .Y(_1167_) );
NAND3X1 NAND3X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(_1167_), .C(_1166_), .Y(_1168_) );
NAND3X1 NAND3X1_216 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(_1164_), .C(_1168_), .Y(_1169_) );
NAND3X1 NAND3X1_217 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf1_), .B(_1167_), .C(_1166_), .Y(_1170_) );
NAND3X1 NAND3X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(_1157_), .C(_1163_), .Y(_1171_) );
NAND3X1 NAND3X1_219 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_1170_), .C(_1171_), .Y(_1172_) );
NAND3X1 NAND3X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1172_), .C(_968_), .Y(_1173_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_746_), .Y(_1174_) );
AOI21X1 AOI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1170_), .B(_1171_), .C(_741_), .Y(_1175_) );
AOI21X1 AOI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1164_), .B(_1168_), .C(_969_), .Y(_1176_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1175_), .B(_1176_), .C(_1174_), .Y(_1177_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_518_), .Y(_1178_) );
NAND3X1 NAND3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1149_), .B(_1150_), .C(_1148_), .Y(_1179_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .B(_1146_), .C(_513_), .Y(_1180_) );
AOI21X1 AOI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1179_), .B(_1180_), .C(bloque_datos_58_bF_buf4_), .Y(_1181_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf3_), .Y(_1182_) );
NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1182_), .B(_1151_), .C(_1147_), .Y(_1183_) );
NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(_1181_), .C(_1183_), .Y(_1184_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1151_), .C(_1182_), .Y(_1185_) );
NAND3X1 NAND3X1_222 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf2_), .B(_1179_), .C(_1180_), .Y(_1186_) );
AOI21X1 AOI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_1185_), .C(_518_), .Y(_1187_) );
NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_1187_), .C(_1184_), .Y(_1188_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_520_), .Y(_1189_) );
NAND3X1 NAND3X1_223 ( .gnd(gnd), .vdd(vdd), .A(_518_), .B(_1186_), .C(_1185_), .Y(_1190_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_1181_), .C(_1178_), .Y(_1191_) );
AOI21X1 AOI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1190_), .B(_1191_), .C(_1189_), .Y(_1192_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1192_), .B(_1188_), .Y(_1193_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_3539_), .B(_3540_), .C(_1193_), .Y(_1194_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_3540_), .B(_3539_), .Y(_1195_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1188_), .B(_1192_), .C(_1195_), .Y(_1196_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1194_), .B(_1196_), .Y(_1197_) );
NAND3X1 NAND3X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1173_), .B(_1197_), .C(_1177_), .Y(_1198_) );
NAND3X1 NAND3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_1164_), .C(_1168_), .Y(_1199_) );
NAND3X1 NAND3X1_226 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(_1170_), .C(_1171_), .Y(_1200_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_759_), .C(_1199_), .D(_1200_), .Y(_1201_) );
AOI21X1 AOI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1172_), .C(_968_), .Y(_1202_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .Y(_1203_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1202_), .B(_1201_), .C(_1203_), .Y(_1204_) );
NAND3X1 NAND3X1_227 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf4_), .B(_1204_), .C(_1198_), .Y(_1205_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf3_), .Y(_1206_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1202_), .B(_1201_), .C(_1197_), .Y(_1207_) );
NAND3X1 NAND3X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1173_), .B(_1203_), .C(_1177_), .Y(_1208_) );
NAND3X1 NAND3X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1206_), .B(_1207_), .C(_1208_), .Y(_1209_) );
NAND3X1 NAND3X1_230 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_1205_), .C(_1209_), .Y(_1210_) );
NAND3X1 NAND3X1_231 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf2_), .B(_1207_), .C(_1208_), .Y(_1211_) );
NAND3X1 NAND3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1206_), .B(_1204_), .C(_1198_), .Y(_1212_) );
NAND3X1 NAND3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_1211_), .C(_1212_), .Y(_1213_) );
NAND3X1 NAND3X1_234 ( .gnd(gnd), .vdd(vdd), .A(_966_), .B(_1210_), .C(_1213_), .Y(_1214_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_966_), .Y(_1215_) );
AOI21X1 AOI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1211_), .B(_1212_), .C(_762_), .Y(_1216_) );
AOI21X1 AOI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(_1209_), .C(_967_), .Y(_1217_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1216_), .B(_1217_), .C(_1215_), .Y(_1218_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf4_), .Y(_1219_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1188_), .B(_1192_), .C(_1219_), .Y(_1220_) );
NAND3X1 NAND3X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1189_), .B(_1190_), .C(_1191_), .Y(_1221_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1184_), .B(_1187_), .C(_521_), .Y(_1222_) );
NAND3X1 NAND3X1_236 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf3_), .B(_1221_), .C(_1222_), .Y(_1223_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1220_), .Y(_1224_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_1224_), .Y(_1225_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_524_), .Y(_1226_) );
AOI21X1 AOI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1220_), .C(_1226_), .Y(_1227_) );
NOR3X1 NOR3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_1227_), .C(_1225_), .Y(_1228_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_525_), .Y(_1229_) );
NAND3X1 NAND3X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .B(_1223_), .C(_1226_), .Y(_1230_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(_1227_), .Y(_1231_) );
AOI21X1 AOI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1230_), .B(_1231_), .C(_1229_), .Y(_1232_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1232_), .B(_1228_), .Y(_1233_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_3551_), .B(_3552_), .C(_1233_), .Y(_1234_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_3552_), .B(_3551_), .Y(_1235_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_1232_), .C(_1235_), .Y(_1236_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1234_), .B(_1236_), .Y(_1237_) );
NAND3X1 NAND3X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1214_), .B(_1237_), .C(_1218_), .Y(_1238_) );
NAND3X1 NAND3X1_239 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_1205_), .C(_1209_), .Y(_1239_) );
NAND3X1 NAND3X1_240 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_1211_), .C(_1212_), .Y(_1240_) );
AOI21X1 AOI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1239_), .B(_1240_), .C(_1215_), .Y(_1241_) );
AOI21X1 AOI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1210_), .B(_1213_), .C(_966_), .Y(_1242_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .Y(_1243_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(_1242_), .C(_1243_), .Y(_1244_) );
NAND3X1 NAND3X1_241 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_134_), .B(_1238_), .C(_1244_), .Y(_1245_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_134_), .Y(_1246_) );
NAND3X1 NAND3X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1214_), .B(_1243_), .C(_1218_), .Y(_1247_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(_1242_), .C(_1237_), .Y(_1248_) );
NAND3X1 NAND3X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1247_), .C(_1248_), .Y(_1249_) );
NAND3X1 NAND3X1_244 ( .gnd(gnd), .vdd(vdd), .A(_964_), .B(_1245_), .C(_1249_), .Y(_1250_) );
NAND3X1 NAND3X1_245 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_134_), .B(_1247_), .C(_1248_), .Y(_1251_) );
NAND3X1 NAND3X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1238_), .C(_1244_), .Y(_1252_) );
NAND3X1 NAND3X1_247 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_1251_), .C(_1252_), .Y(_1253_) );
NAND3X1 NAND3X1_248 ( .gnd(gnd), .vdd(vdd), .A(_963_), .B(_1250_), .C(_1253_), .Y(_1254_) );
INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(_963_), .Y(_1255_) );
AOI21X1 AOI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1251_), .B(_1252_), .C(_789_), .Y(_1256_) );
AOI21X1 AOI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1245_), .B(_1249_), .C(_964_), .Y(_1257_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_1257_), .C(_1255_), .Y(_1258_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_530_), .Y(_1259_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf4_), .Y(_1260_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_1232_), .C(_1260_), .Y(_1261_) );
NAND3X1 NAND3X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1229_), .B(_1230_), .C(_1231_), .Y(_1262_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .B(_1227_), .C(_527_), .Y(_1263_) );
NAND3X1 NAND3X1_250 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf3_), .B(_1263_), .C(_1262_), .Y(_1264_) );
NAND3X1 NAND3X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .B(_1264_), .C(_1259_), .Y(_1265_) );
AOI21X1 AOI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1263_), .B(_1262_), .C(bloque_datos_90_bF_buf2_), .Y(_1266_) );
NOR3X1 NOR3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1232_), .B(_1260_), .C(_1228_), .Y(_1267_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1266_), .C(_530_), .Y(_1268_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .B(_1265_), .Y(_1269_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_1269_), .Y(_1270_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_1270_), .Y(_1271_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_1269_), .Y(_1272_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .B(_1271_), .Y(_1273_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(_1273_), .Y(_1274_) );
NAND3X1 NAND3X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1254_), .B(_1274_), .C(_1258_), .Y(_1275_) );
NAND3X1 NAND3X1_253 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_1245_), .C(_1249_), .Y(_1276_) );
NAND3X1 NAND3X1_254 ( .gnd(gnd), .vdd(vdd), .A(_964_), .B(_1251_), .C(_1252_), .Y(_1277_) );
AOI21X1 AOI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_1277_), .C(_1255_), .Y(_1278_) );
AOI21X1 AOI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1250_), .B(_1253_), .C(_963_), .Y(_1279_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .B(_1279_), .C(_1273_), .Y(_1280_) );
NAND3X1 NAND3X1_255 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_1275_), .C(_1280_), .Y(_1281_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_150_), .B(_1281_), .Y(_1282_) );
INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_150_), .Y(_1283_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .B(_1279_), .C(_1274_), .Y(_1284_) );
NAND3X1 NAND3X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1254_), .B(_1273_), .C(_1258_), .Y(_1285_) );
AOI21X1 AOI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1285_), .B(_1284_), .C(_961_), .Y(_1286_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(_1286_), .Y(_1287_) );
NAND3X1 NAND3X1_257 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_1282_), .C(_1287_), .Y(_1288_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_150_), .B(_1286_), .Y(_1289_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(_1281_), .Y(_1290_) );
NAND3X1 NAND3X1_258 ( .gnd(gnd), .vdd(vdd), .A(_806_), .B(_1290_), .C(_1289_), .Y(_1291_) );
AOI21X1 AOI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1288_), .B(_1291_), .C(_960_), .Y(_1292_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_818_), .Y(_1293_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1293_), .B(_610_), .C(_817_), .Y(_1294_) );
NAND3X1 NAND3X1_259 ( .gnd(gnd), .vdd(vdd), .A(_806_), .B(_1282_), .C(_1287_), .Y(_1295_) );
NAND3X1 NAND3X1_260 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_1290_), .C(_1289_), .Y(_1296_) );
AOI21X1 AOI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1296_), .C(_1294_), .Y(_1297_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_138_), .Y(_1298_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1271_), .B(_1272_), .C(_1298_), .Y(_1299_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_138_), .B(_1273_), .Y(_1300_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_1300_), .Y(_1301_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_1301_), .Y(_1302_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_1302_), .Y(_1303_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_535_), .C(_1301_), .Y(_1304_) );
NAND3X1 NAND3X1_261 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_1304_), .C(_1303_), .Y(_1305_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(_1304_), .Y(_1306_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_1302_), .C(_542_), .Y(_1307_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(_1305_), .Y(_1308_) );
INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(_1308_), .Y(_1309_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_1297_), .C(_1309_), .Y(_1310_) );
NAND3X1 NAND3X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1296_), .C(_1294_), .Y(_1311_) );
AOI21X1 AOI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .B(_1289_), .C(_812_), .Y(_1312_) );
AOI21X1 AOI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1282_), .B(_1287_), .C(_806_), .Y(_1313_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(_1313_), .C(_960_), .Y(_1314_) );
NAND3X1 NAND3X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1308_), .B(_1311_), .C(_1314_), .Y(_1315_) );
NAND3X1 NAND3X1_264 ( .gnd(gnd), .vdd(vdd), .A(_3787_), .B(_1315_), .C(_1310_), .Y(_1316_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_166_), .B(_1316_), .Y(_1317_) );
INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_166_), .Y(_1318_) );
NAND3X1 NAND3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(_1311_), .C(_1314_), .Y(_1319_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_1297_), .C(_1308_), .Y(_1320_) );
AOI21X1 AOI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1319_), .B(_1320_), .C(_3574_), .Y(_1321_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1318_), .B(_1321_), .Y(_1322_) );
NAND3X1 NAND3X1_266 ( .gnd(gnd), .vdd(vdd), .A(_831_), .B(_1317_), .C(_1322_), .Y(_1323_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_166_), .B(_1321_), .Y(_1324_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1318_), .B(_1316_), .Y(_1325_) );
NAND3X1 NAND3X1_267 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_1325_), .C(_1324_), .Y(_1326_) );
AOI21X1 AOI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1323_), .B(_1326_), .C(_958_), .Y(_1327_) );
NOR3X1 NOR3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(_607_), .C(_831_), .Y(_1328_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1328_), .B(_606_), .C(_836_), .Y(_1329_) );
NAND3X1 NAND3X1_268 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_1317_), .C(_1322_), .Y(_1330_) );
NAND3X1 NAND3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_831_), .B(_1325_), .C(_1324_), .Y(_1331_) );
AOI21X1 AOI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1330_), .B(_1331_), .C(_1329_), .Y(_1332_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_154_), .Y(_1333_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .B(_1308_), .Y(_1334_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .B(_1308_), .Y(_1335_) );
INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(_1335_), .Y(_1336_) );
NAND3X1 NAND3X1_270 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_1334_), .C(_1336_), .Y(_1337_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_1334_), .Y(_1338_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .B(_1335_), .C(_546_), .Y(_1339_) );
NAND3X1 NAND3X1_271 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_1339_), .C(_1337_), .Y(_1340_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1339_), .B(_1337_), .Y(_1341_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_547_), .C(_1341_), .Y(_1342_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(_1342_), .Y(_1343_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .Y(_1344_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1327_), .B(_1332_), .C(_1344_), .Y(_1345_) );
NAND3X1 NAND3X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1329_), .B(_1330_), .C(_1331_), .Y(_1346_) );
AOI21X1 AOI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1325_), .B(_1324_), .C(_831_), .Y(_1347_) );
AOI21X1 AOI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1322_), .C(_825_), .Y(_1348_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1347_), .B(_1348_), .C(_958_), .Y(_1349_) );
NAND3X1 NAND3X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_1346_), .C(_1349_), .Y(_1350_) );
NAND3X1 NAND3X1_274 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_1350_), .C(_1345_), .Y(_1351_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_182_), .B(_1351_), .Y(_1352_) );
INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_182_), .Y(_1353_) );
NAND3X1 NAND3X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1344_), .B(_1346_), .C(_1349_), .Y(_1354_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1327_), .B(_1332_), .C(_1343_), .Y(_1355_) );
AOI21X1 AOI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1354_), .B(_1355_), .C(_3584_), .Y(_1356_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1353_), .B(_1356_), .Y(_1357_) );
NAND3X1 NAND3X1_276 ( .gnd(gnd), .vdd(vdd), .A(_842_), .B(_1352_), .C(_1357_), .Y(_1358_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1354_), .B(_1355_), .Y(_1359_) );
NAND3X1 NAND3X1_277 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_182_), .B(_956_), .C(_1359_), .Y(_1360_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1353_), .B(_1351_), .Y(_1361_) );
NAND3X1 NAND3X1_278 ( .gnd(gnd), .vdd(vdd), .A(_849_), .B(_1360_), .C(_1361_), .Y(_1362_) );
NAND3X1 NAND3X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1362_), .B(_955_), .C(_1358_), .Y(_1363_) );
AOI21X1 AOI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_842_), .B(_847_), .C(_352_), .Y(_1364_) );
AOI21X1 AOI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_853_), .C(_1364_), .Y(_1365_) );
AOI21X1 AOI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_1361_), .C(_849_), .Y(_1366_) );
AOI21X1 AOI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .B(_1357_), .C(_842_), .Y(_1367_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1367_), .B(_1366_), .C(_1365_), .Y(_1368_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(_558_), .Y(_1369_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_170_), .Y(_1370_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1370_), .B(_1343_), .Y(_1371_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_1371_), .Y(_1372_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1370_), .B(_1343_), .Y(_1373_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .B(_1372_), .Y(_1374_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .B(_555_), .Y(_1375_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .B(_1373_), .C(_554_), .Y(_1376_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_1376_), .Y(_1377_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1377_), .B(_1375_), .Y(_1378_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1369_), .B(_1378_), .Y(_1379_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1375_), .B(_1377_), .C(_558_), .Y(_1380_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1380_), .B(_1379_), .Y(_1381_) );
NAND3X1 NAND3X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_1381_), .C(_1368_), .Y(_1382_) );
NAND3X1 NAND3X1_281 ( .gnd(gnd), .vdd(vdd), .A(_849_), .B(_1352_), .C(_1357_), .Y(_1383_) );
NAND3X1 NAND3X1_282 ( .gnd(gnd), .vdd(vdd), .A(_842_), .B(_1360_), .C(_1361_), .Y(_1384_) );
AOI21X1 AOI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1384_), .B(_1383_), .C(_1365_), .Y(_1385_) );
AOI21X1 AOI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1362_), .B(_1358_), .C(_955_), .Y(_1386_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_1381_), .Y(_1387_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1385_), .B(_1386_), .C(_1387_), .Y(_1388_) );
NAND3X1 NAND3X1_283 ( .gnd(gnd), .vdd(vdd), .A(_953_), .B(_1382_), .C(_1388_), .Y(_1389_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_198_), .B(_1389_), .Y(_1390_) );
INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_198_), .Y(_1391_) );
AOI21X1 AOI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_1368_), .C(_1381_), .Y(_1392_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_1392_), .Y(_1393_) );
NAND3X1 NAND3X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1391_), .B(_1382_), .C(_1393_), .Y(_1394_) );
NAND3X1 NAND3X1_285 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_1390_), .C(_1394_), .Y(_1395_) );
NAND3X1 NAND3X1_286 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_198_), .B(_1382_), .C(_1393_), .Y(_1396_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1391_), .B(_1389_), .Y(_1397_) );
NAND3X1 NAND3X1_287 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_1397_), .C(_1396_), .Y(_1398_) );
AOI21X1 AOI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_1398_), .C(_951_), .Y(_1399_) );
NOR3X1 NOR3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_601_), .C(_868_), .Y(_1400_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1400_), .B(_600_), .C(_873_), .Y(_1401_) );
NAND3X1 NAND3X1_288 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_1390_), .C(_1394_), .Y(_1402_) );
NAND3X1 NAND3X1_289 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_1397_), .C(_1396_), .Y(_1403_) );
AOI21X1 AOI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1402_), .B(_1403_), .C(_1401_), .Y(_1404_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_566_), .Y(_1405_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_186_), .Y(_1406_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1406_), .B(_1381_), .Y(_1407_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1406_), .B(_1381_), .Y(_1408_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .Y(_1409_) );
NAND3X1 NAND3X1_290 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_1407_), .C(_1409_), .Y(_1410_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(_1407_), .Y(_1411_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1411_), .B(_1408_), .C(_562_), .Y(_1412_) );
NAND3X1 NAND3X1_291 ( .gnd(gnd), .vdd(vdd), .A(_1405_), .B(_1412_), .C(_1410_), .Y(_1413_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(_1410_), .Y(_1414_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_1412_), .Y(_1415_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(_1415_), .C(_566_), .Y(_1416_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1413_), .B(_1416_), .Y(_1417_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .Y(_1418_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1399_), .B(_1404_), .C(_1418_), .Y(_1419_) );
NAND3X1 NAND3X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1402_), .B(_1403_), .C(_1401_), .Y(_1420_) );
AOI21X1 AOI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1397_), .B(_1396_), .C(_868_), .Y(_1421_) );
AOI21X1 AOI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1390_), .B(_1394_), .C(_862_), .Y(_1422_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1421_), .B(_1422_), .C(_951_), .Y(_1423_) );
NAND3X1 NAND3X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1417_), .C(_1423_), .Y(_1424_) );
NAND3X1 NAND3X1_294 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(_1424_), .C(_1419_), .Y(_1425_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_214_), .B(_1425_), .Y(_1426_) );
INVX2 INVX2_42 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_214_), .Y(_1427_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1399_), .B(_1404_), .C(_1417_), .Y(_1428_) );
NAND3X1 NAND3X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1418_), .C(_1423_), .Y(_1429_) );
AOI21X1 AOI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1429_), .B(_1428_), .C(_3602_), .Y(_1430_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1427_), .B(_1430_), .Y(_1431_) );
NAND3X1 NAND3X1_296 ( .gnd(gnd), .vdd(vdd), .A(_887_), .B(_1426_), .C(_1431_), .Y(_1432_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_214_), .B(_1430_), .Y(_1433_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1427_), .B(_1425_), .Y(_1434_) );
NAND3X1 NAND3X1_297 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_1434_), .C(_1433_), .Y(_1435_) );
AOI21X1 AOI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1432_), .B(_1435_), .C(_948_), .Y(_1436_) );
NOR3X1 NOR3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_888_), .B(_598_), .C(_887_), .Y(_1437_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1437_), .B(_597_), .C(_892_), .Y(_1438_) );
NAND3X1 NAND3X1_298 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_1426_), .C(_1431_), .Y(_1439_) );
NAND3X1 NAND3X1_299 ( .gnd(gnd), .vdd(vdd), .A(_887_), .B(_1434_), .C(_1433_), .Y(_1440_) );
AOI21X1 AOI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(_1440_), .C(_1438_), .Y(_1441_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_574_), .Y(_1442_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_202_), .Y(_1443_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1443_), .B(_1417_), .Y(_1444_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1443_), .B(_1417_), .Y(_1445_) );
INVX2 INVX2_43 ( .gnd(gnd), .vdd(vdd), .A(_1445_), .Y(_1446_) );
NAND3X1 NAND3X1_300 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_1444_), .C(_1446_), .Y(_1447_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(_1444_), .Y(_1448_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1448_), .B(_1445_), .C(_570_), .Y(_1449_) );
NAND3X1 NAND3X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1442_), .B(_1449_), .C(_1447_), .Y(_1450_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .Y(_1451_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_1449_), .Y(_1452_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1451_), .B(_1452_), .C(_574_), .Y(_1453_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .B(_1453_), .Y(_1454_) );
INVX2 INVX2_44 ( .gnd(gnd), .vdd(vdd), .A(_1454_), .Y(_1455_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1441_), .B(_1436_), .C(_1455_), .Y(_1456_) );
NAND3X1 NAND3X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(_1440_), .C(_1438_), .Y(_1457_) );
AOI21X1 AOI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_1433_), .C(_887_), .Y(_1458_) );
AOI21X1 AOI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(_1431_), .C(_881_), .Y(_1459_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1458_), .B(_1459_), .C(_948_), .Y(_1460_) );
NAND3X1 NAND3X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1454_), .B(_1460_), .C(_1457_), .Y(_1461_) );
NAND3X1 NAND3X1_304 ( .gnd(gnd), .vdd(vdd), .A(_946_), .B(_1461_), .C(_1456_), .Y(_1462_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_230_), .B(_1462_), .Y(_1463_) );
INVX2 INVX2_45 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_230_), .Y(_1464_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1441_), .B(_1436_), .C(_1454_), .Y(_1465_) );
NAND3X1 NAND3X1_305 ( .gnd(gnd), .vdd(vdd), .A(_1455_), .B(_1460_), .C(_1457_), .Y(_1466_) );
AOI21X1 AOI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_1465_), .C(_945_), .Y(_1467_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_1467_), .Y(_1468_) );
NAND3X1 NAND3X1_306 ( .gnd(gnd), .vdd(vdd), .A(_906_), .B(_1463_), .C(_1468_), .Y(_1469_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_230_), .B(_1467_), .Y(_1470_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_1462_), .Y(_1471_) );
NAND3X1 NAND3X1_307 ( .gnd(gnd), .vdd(vdd), .A(_900_), .B(_1471_), .C(_1470_), .Y(_1472_) );
AOI21X1 AOI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(_1472_), .C(_942_), .Y(_1473_) );
NOR3X1 NOR3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_907_), .B(_595_), .C(_906_), .Y(_1474_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1474_), .B(_594_), .C(_911_), .Y(_1475_) );
NAND3X1 NAND3X1_308 ( .gnd(gnd), .vdd(vdd), .A(_900_), .B(_1463_), .C(_1468_), .Y(_1476_) );
NAND3X1 NAND3X1_309 ( .gnd(gnd), .vdd(vdd), .A(_906_), .B(_1471_), .C(_1470_), .Y(_1477_) );
AOI21X1 AOI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1476_), .B(_1477_), .C(_1475_), .Y(_1478_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(_582_), .Y(_1479_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_218_), .Y(_1480_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1480_), .B(_1454_), .Y(_1481_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1480_), .B(_1454_), .Y(_1482_) );
INVX2 INVX2_46 ( .gnd(gnd), .vdd(vdd), .A(_1482_), .Y(_1483_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1481_), .B(_1483_), .Y(_1484_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .B(_578_), .Y(_1485_) );
AOI21X1 AOI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1481_), .B(_1483_), .C(_579_), .Y(_1486_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(_1486_), .Y(_1487_) );
NAND3X1 NAND3X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1479_), .B(_1487_), .C(_1485_), .Y(_1488_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_578_), .B(_1484_), .Y(_1489_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1489_), .B(_1486_), .C(_582_), .Y(_1490_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1490_), .B(_1488_), .Y(_1491_) );
INVX2 INVX2_47 ( .gnd(gnd), .vdd(vdd), .A(_1491_), .Y(_1492_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1478_), .B(_1473_), .C(_1492_), .Y(_1493_) );
NAND3X1 NAND3X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1476_), .B(_1477_), .C(_1475_), .Y(_1494_) );
AOI21X1 AOI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .B(_1470_), .C(_906_), .Y(_1495_) );
AOI21X1 AOI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_1468_), .C(_900_), .Y(_1496_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1495_), .B(_1496_), .C(_942_), .Y(_1497_) );
NAND3X1 NAND3X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1497_), .B(_1491_), .C(_1494_), .Y(_1498_) );
NAND3X1 NAND3X1_313 ( .gnd(gnd), .vdd(vdd), .A(_3852_), .B(_1498_), .C(_1493_), .Y(_1499_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_246_), .B(_1499_), .Y(_1500_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_246_), .Y(_1501_) );
NAND3X1 NAND3X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1497_), .B(_1492_), .C(_1494_), .Y(_1502_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1478_), .B(_1473_), .C(_1491_), .Y(_1503_) );
AOI21X1 AOI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_1503_), .C(_3624_), .Y(_1504_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1501_), .B(_1504_), .Y(_1505_) );
NAND3X1 NAND3X1_315 ( .gnd(gnd), .vdd(vdd), .A(_925_), .B(_1500_), .C(_1505_), .Y(_1506_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_246_), .B(_1504_), .Y(_1507_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1501_), .B(_1499_), .Y(_1508_) );
NAND3X1 NAND3X1_316 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_1508_), .C(_1507_), .Y(_1509_) );
AOI21X1 AOI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .B(_1509_), .C(_940_), .Y(_1510_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_929_), .C(_927_), .Y(_1511_) );
NAND3X1 NAND3X1_317 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_1500_), .C(_1505_), .Y(_1512_) );
NAND3X1 NAND3X1_318 ( .gnd(gnd), .vdd(vdd), .A(_925_), .B(_1508_), .C(_1507_), .Y(_1513_) );
AOI21X1 AOI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1512_), .B(_1513_), .C(_1511_), .Y(_1514_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(_590_), .Y(_1515_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_234_), .B(_1492_), .Y(_1516_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(_1516_), .Y(_1517_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_234_), .B(_1492_), .Y(_1518_) );
NAND3X1 NAND3X1_319 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_1518_), .C(_1517_), .Y(_1519_) );
INVX2 INVX2_48 ( .gnd(gnd), .vdd(vdd), .A(_1518_), .Y(_1520_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1520_), .B(_1516_), .C(_586_), .Y(_1521_) );
NAND3X1 NAND3X1_320 ( .gnd(gnd), .vdd(vdd), .A(_1515_), .B(_1521_), .C(_1519_), .Y(_1522_) );
NOR3X1 NOR3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_1516_), .C(_1520_), .Y(_1523_) );
AOI21X1 AOI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1518_), .B(_1517_), .C(_587_), .Y(_1524_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1523_), .C(_590_), .Y(_1525_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1522_), .B(_1525_), .Y(_1526_) );
INVX2 INVX2_49 ( .gnd(gnd), .vdd(vdd), .A(_1526_), .Y(_1527_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1514_), .B(_1510_), .C(_1527_), .Y(_1528_) );
NAND3X1 NAND3X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1512_), .B(_1513_), .C(_1511_), .Y(_1529_) );
NAND3X1 NAND3X1_322 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .B(_1509_), .C(_940_), .Y(_1530_) );
NAND3X1 NAND3X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1530_), .B(_1526_), .C(_1529_), .Y(_1531_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1531_), .B(_1528_), .Y(_1532_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_939_), .Y(module_0_H_6_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1514_), .B(_1510_), .C(_1526_), .Y(_1533_) );
NAND3X1 NAND3X1_324 ( .gnd(gnd), .vdd(vdd), .A(_1530_), .B(_1527_), .C(_1529_), .Y(_1534_) );
NAND3X1 NAND3X1_325 ( .gnd(gnd), .vdd(vdd), .A(_1534_), .B(_1533_), .C(_939_), .Y(_1535_) );
AOI21X1 AOI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1508_), .B(_1507_), .C(_925_), .Y(_1536_) );
AOI21X1 AOI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1513_), .B(_1511_), .C(_1536_), .Y(_1537_) );
AOI21X1 AOI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1515_), .B(_1521_), .C(_1523_), .Y(_1538_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_1486_), .C(_1485_), .Y(_1539_) );
AOI21X1 AOI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1442_), .B(_1449_), .C(_1451_), .Y(_1540_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_203_), .Y(_1541_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1415_), .B(_566_), .C(_1410_), .Y(_1542_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_187_), .Y(_1543_) );
AOI21X1 AOI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1369_), .B(_1376_), .C(_1375_), .Y(_1544_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .Y(_1545_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .Y(_1546_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_171_), .Y(_1547_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .B(_550_), .C(_1337_), .Y(_1548_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_155_), .Y(_1549_) );
AOI21X1 AOI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_1304_), .C(_1302_), .Y(_1550_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .Y(_1551_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1551_), .B(_534_), .C(_1265_), .Y(_1552_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_1227_), .C(_1230_), .Y(_1553_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .Y(_1554_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_1187_), .C(_1190_), .Y(_1555_) );
AOI21X1 AOI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1148_), .B(_1150_), .C(_1143_), .Y(_1556_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf3_), .Y(_1557_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_504_), .Y(_1558_) );
AOI21X1 AOI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1558_), .B(_1107_), .C(_1110_), .Y(_1559_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(_1071_), .Y(_1560_) );
AOI21X1 AOI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1064_), .B(_1560_), .C(_1070_), .Y(_1561_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .Y(_1562_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .Y(_1563_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1038_), .B(_1035_), .C(_1031_), .Y(_1564_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_27_), .B(module_0_W_11_), .Y(_1565_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(_1565_), .Y(_1566_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_27_), .B(module_0_W_11_), .Y(_1567_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1567_), .B(_1566_), .Y(_1568_) );
NAND3X1 NAND3X1_326 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_26_), .B(module_0_W_10_), .C(_1568_), .Y(_1569_) );
NAND3X1 NAND3X1_327 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .B(_1567_), .C(_1566_), .Y(_1570_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1570_), .B(_1569_), .Y(_1571_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1564_), .B(_1571_), .Y(_1572_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1563_), .B(_1572_), .Y(_1573_) );
XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1564_), .B(_1571_), .Y(_1574_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .B(_1574_), .Y(_1575_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1575_), .B(_1573_), .Y(_1576_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .B(_1576_), .Y(_1577_) );
NAND3X1 NAND3X1_328 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1575_), .C(_1573_), .Y(_1578_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1578_), .B(_1577_), .Y(_1579_) );
XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1579_), .B(_1561_), .Y(_1580_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf4_), .B(_1580_), .Y(_1581_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf3_), .Y(_1582_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .B(_1065_), .Y(_1583_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_1071_), .C(_1583_), .Y(_1584_) );
XNOR2X1 XNOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1579_), .B(_1584_), .Y(_1585_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .B(_1585_), .Y(_1586_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1581_), .B(_1586_), .Y(_1587_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1587_), .Y(_1588_) );
AOI21X1 AOI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1581_), .B(_1586_), .C(_1106_), .Y(_1589_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1588_), .B(_1589_), .C(_1559_), .Y(_1590_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1111_), .B(_505_), .C(_1103_), .Y(_1591_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .B(_1102_), .Y(_1592_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(_1589_), .Y(_1593_) );
NAND3X1 NAND3X1_329 ( .gnd(gnd), .vdd(vdd), .A(_1593_), .B(_1591_), .C(_1592_), .Y(_1594_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1590_), .B(_1594_), .Y(_1595_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1557_), .B(_1595_), .Y(_1596_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_1594_), .B(_1590_), .Y(_1597_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf2_), .B(_1597_), .Y(_1598_) );
AOI21X1 AOI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1596_), .B(_1598_), .C(_1145_), .Y(_1599_) );
NAND3X1 NAND3X1_330 ( .gnd(gnd), .vdd(vdd), .A(_1145_), .B(_1596_), .C(_1598_), .Y(_1600_) );
INVX2 INVX2_50 ( .gnd(gnd), .vdd(vdd), .A(_1600_), .Y(_1601_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1601_), .B(_1599_), .C(_1556_), .Y(_1602_) );
INVX2 INVX2_51 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .Y(_1603_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1599_), .B(_1601_), .Y(_1604_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .B(_1147_), .C(_1604_), .Y(_1605_) );
INVX2 INVX2_52 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .Y(_1606_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .B(_1603_), .C(bloque_datos_59_bF_buf4_), .Y(_1607_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf3_), .Y(_1608_) );
NAND3X1 NAND3X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .B(_1602_), .C(_1605_), .Y(_1609_) );
NAND3X1 NAND3X1_332 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_1609_), .C(_1607_), .Y(_1610_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .B(_1603_), .C(_1608_), .Y(_1611_) );
NAND3X1 NAND3X1_333 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf2_), .B(_1602_), .C(_1605_), .Y(_1612_) );
NAND3X1 NAND3X1_334 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_1612_), .C(_1611_), .Y(_1613_) );
AOI21X1 AOI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1610_), .B(_1613_), .C(_1555_), .Y(_1614_) );
NAND3X1 NAND3X1_335 ( .gnd(gnd), .vdd(vdd), .A(_1555_), .B(_1610_), .C(_1613_), .Y(_1615_) );
INVX2 INVX2_53 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .Y(_1616_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1616_), .B(_1614_), .C(bloque_datos_75_bF_buf4_), .Y(_1617_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf3_), .Y(_1618_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(_1614_), .Y(_1619_) );
NAND3X1 NAND3X1_336 ( .gnd(gnd), .vdd(vdd), .A(_1618_), .B(_1615_), .C(_1619_), .Y(_1620_) );
NAND3X1 NAND3X1_337 ( .gnd(gnd), .vdd(vdd), .A(_1554_), .B(_1620_), .C(_1617_), .Y(_1621_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1616_), .B(_1614_), .C(_1618_), .Y(_1622_) );
NAND3X1 NAND3X1_338 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf2_), .B(_1615_), .C(_1619_), .Y(_1623_) );
NAND3X1 NAND3X1_339 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1623_), .C(_1622_), .Y(_1624_) );
AOI21X1 AOI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(_1624_), .C(_1553_), .Y(_1625_) );
NAND3X1 NAND3X1_340 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1621_), .C(_1624_), .Y(_1626_) );
INVX2 INVX2_54 ( .gnd(gnd), .vdd(vdd), .A(_1626_), .Y(_1627_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .B(_1625_), .C(bloque_datos_91_bF_buf3_), .Y(_1628_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf2_), .Y(_1629_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .Y(_1630_) );
NAND3X1 NAND3X1_341 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(_1626_), .C(_1630_), .Y(_1631_) );
NAND3X1 NAND3X1_342 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1631_), .C(_1628_), .Y(_1632_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .B(_1625_), .C(_1629_), .Y(_1633_) );
NAND3X1 NAND3X1_343 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf1_), .B(_1626_), .C(_1630_), .Y(_1634_) );
NAND3X1 NAND3X1_344 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .B(_1634_), .C(_1633_), .Y(_1635_) );
NAND3X1 NAND3X1_345 ( .gnd(gnd), .vdd(vdd), .A(_1632_), .B(_1635_), .C(_1552_), .Y(_1636_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .Y(_1637_) );
AOI21X1 AOI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1632_), .B(_1635_), .C(_1552_), .Y(_1638_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1638_), .B(_1637_), .Y(_1639_) );
XNOR2X1 XNOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(module_0_W_139_), .Y(_1640_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1300_), .B(_1640_), .Y(_1641_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .Y(_1642_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1298_), .B(_1274_), .C(_1640_), .Y(_1643_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(_1642_), .Y(_1644_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_1644_), .B(_1550_), .Y(_1645_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .Y(_1646_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1646_), .B(_1641_), .C(_1550_), .Y(_1647_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(_1645_), .Y(_1648_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1549_), .B(_1648_), .Y(_1649_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .Y(_1650_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1549_), .B(_1648_), .Y(_1651_) );
NOR3X1 NOR3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1651_), .C(_1650_), .Y(_1652_) );
INVX2 INVX2_55 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .Y(_1653_) );
AOI21X1 AOI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .B(_1653_), .C(_1335_), .Y(_1654_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1652_), .B(_1654_), .Y(_1655_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1548_), .Y(_1656_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(_1337_), .Y(_1657_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1654_), .B(_1652_), .C(_1657_), .Y(_1658_) );
INVX2 INVX2_56 ( .gnd(gnd), .vdd(vdd), .A(_1658_), .Y(_1659_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1656_), .B(_1659_), .C(_1547_), .Y(_1660_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1659_), .B(_1656_), .Y(_1661_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_171_), .B(_1661_), .Y(_1662_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1662_), .Y(_1663_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1546_), .B(_1663_), .Y(_1664_) );
AOI21X1 AOI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1662_), .C(_1373_), .Y(_1665_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .B(_1664_), .Y(_1666_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_1666_), .B(_1545_), .Y(_1667_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1664_), .B(_1665_), .C(_1544_), .Y(_1668_) );
INVX2 INVX2_57 ( .gnd(gnd), .vdd(vdd), .A(_1668_), .Y(_1669_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1667_), .B(_1669_), .C(_1543_), .Y(_1670_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1669_), .B(_1667_), .Y(_1671_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_187_), .B(_1671_), .Y(_1672_) );
NAND3X1 NAND3X1_346 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .B(_1670_), .C(_1672_), .Y(_1673_) );
INVX2 INVX2_58 ( .gnd(gnd), .vdd(vdd), .A(_1673_), .Y(_1674_) );
AOI21X1 AOI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1670_), .B(_1672_), .C(_1408_), .Y(_1675_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1675_), .B(_1674_), .Y(_1676_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1542_), .B(_1676_), .Y(_1677_) );
AOI21X1 AOI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1405_), .B(_1412_), .C(_1414_), .Y(_1678_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1674_), .B(_1675_), .C(_1678_), .Y(_1679_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1679_), .B(_1677_), .Y(_1680_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(_1680_), .Y(_1681_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(_1680_), .Y(_1682_) );
INVX2 INVX2_59 ( .gnd(gnd), .vdd(vdd), .A(_1682_), .Y(_1683_) );
NAND3X1 NAND3X1_347 ( .gnd(gnd), .vdd(vdd), .A(_1445_), .B(_1681_), .C(_1683_), .Y(_1684_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .Y(_1685_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1685_), .B(_1682_), .C(_1446_), .Y(_1686_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1686_), .B(_1684_), .Y(_1687_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1540_), .B(_1687_), .Y(_1688_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1452_), .B(_574_), .C(_1447_), .Y(_1689_) );
AOI21X1 AOI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1686_), .B(_1684_), .C(_1689_), .Y(_1690_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1690_), .B(_1688_), .Y(_1691_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_219_), .B(_1691_), .Y(_1692_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_1691_), .B(module_0_W_219_), .Y(_1693_) );
NOR3X1 NOR3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_1483_), .C(_1693_), .Y(_1694_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_1691_), .B(module_0_W_219_), .Y(_1695_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_219_), .B(_1691_), .Y(_1696_) );
AOI21X1 AOI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1696_), .B(_1695_), .C(_1482_), .Y(_1697_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(_1694_), .Y(_1698_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_1698_), .B(_1539_), .Y(_1699_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1539_), .B(_1698_), .Y(_1700_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1700_), .B(_1699_), .Y(_1701_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_1701_), .B(module_0_W_235_), .Y(_1702_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_235_), .B(_1701_), .Y(_1703_) );
NAND3X1 NAND3X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1520_), .B(_1703_), .C(_1702_), .Y(_1704_) );
INVX2 INVX2_60 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .Y(_1705_) );
AOI21X1 AOI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1703_), .B(_1702_), .C(_1520_), .Y(_1706_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .B(_1706_), .C(_1538_), .Y(_1707_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(_1707_), .Y(_1708_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_590_), .C(_1519_), .Y(_1709_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1706_), .B(_1705_), .Y(_1710_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_1710_), .B(_1709_), .Y(_1711_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1708_), .B(_1711_), .Y(_1712_) );
INVX2 INVX2_61 ( .gnd(gnd), .vdd(vdd), .A(_1712_), .Y(_1713_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(_1701_), .Y(_1714_) );
AOI21X1 AOI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1403_), .B(_1401_), .C(_1421_), .Y(_1715_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1367_), .B(_1365_), .C(_1358_), .Y(_1716_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(_1716_), .Y(_1717_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_1667_), .B(_1669_), .Y(_1718_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1321_), .B(_1318_), .C(module_0_W_167_), .Y(_1719_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_167_), .Y(_1720_) );
NAND3X1 NAND3X1_349 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_166_), .B(_1720_), .C(_1316_), .Y(_1721_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_1656_), .B(_1659_), .Y(_1722_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(_1245_), .Y(_1723_) );
AOI21X1 AOI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_966_), .B(_1213_), .C(_1216_), .Y(_1724_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .Y(_1725_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .B(_1627_), .Y(_1726_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_1176_), .C(_1169_), .Y(_1727_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1614_), .B(_1616_), .Y(_1728_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .B(_1134_), .C(_1127_), .Y(_1729_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1603_), .B(_1606_), .Y(_1730_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(_1730_), .Y(_1731_) );
AOI21X1 AOI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1092_), .B(_972_), .C(_1095_), .Y(_1732_) );
AOI21X1 AOI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_974_), .C(_1060_), .Y(_1733_) );
AOI21X1 AOI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_977_), .B(_1019_), .C(_1023_), .Y(_1734_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(_994_), .Y(_1735_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .B(_999_), .Y(_1736_) );
XNOR2X1 XNOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_7_), .B(module_0_W_23_), .Y(_1737_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .B(_1737_), .Y(_1738_) );
XNOR2X1 XNOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_985_), .B(module_0_W_11_), .Y(_1739_) );
XNOR2X1 XNOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1739_), .B(_1738_), .Y(_1740_) );
XNOR2X1 XNOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1740_), .B(_989_), .Y(_1741_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_3683_), .B(_3685_), .Y(_1742_) );
XNOR2X1 XNOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1742_), .B(bloque_datos[7]), .Y(_1743_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1741_), .B(_1743_), .Y(_1744_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_1743_), .B(_1741_), .Y(_1745_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1744_), .B(_1745_), .Y(_1746_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .B(_1746_), .Y(_1747_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .B(_1736_), .Y(_1748_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1748_), .B(_1747_), .C(_1572_), .Y(_1749_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .B(_1736_), .Y(_1750_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .B(_1746_), .Y(_1751_) );
NAND3X1 NAND3X1_350 ( .gnd(gnd), .vdd(vdd), .A(_1574_), .B(_1751_), .C(_1750_), .Y(_1752_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_1752_), .B(_1749_), .Y(_1753_) );
AOI21X1 AOI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_1013_), .C(_1012_), .Y(_1754_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_3702_), .B(_3697_), .C(bloque_datos_23_bF_buf3_), .Y(_1755_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(_3698_), .Y(_1756_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_1756_), .B(bloque_datos_23_bF_buf2_), .Y(_1757_) );
NAND3X1 NAND3X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1755_), .B(_1754_), .C(_1757_), .Y(_1758_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(_1755_), .Y(_1759_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf1_), .B(_1756_), .Y(_1760_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1760_), .B(_1759_), .C(_1011_), .Y(_1761_) );
AOI21X1 AOI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1758_), .B(_1761_), .C(_1753_), .Y(_1762_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1749_), .B(_1752_), .Y(_1763_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1761_), .B(_1758_), .Y(_1764_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1763_), .B(_1764_), .Y(_1765_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1765_), .B(_1762_), .C(_1734_), .Y(_1766_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(_1734_), .Y(_1767_) );
NOR3X1 NOR3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1760_), .B(_1759_), .C(_1011_), .Y(_1768_) );
AOI21X1 AOI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1755_), .B(_1757_), .C(_1754_), .Y(_1769_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1768_), .B(_1769_), .C(_1763_), .Y(_1770_) );
NAND3X1 NAND3X1_352 ( .gnd(gnd), .vdd(vdd), .A(_1758_), .B(_1761_), .C(_1753_), .Y(_1771_) );
NAND3X1 NAND3X1_353 ( .gnd(gnd), .vdd(vdd), .A(_1770_), .B(_1771_), .C(_1767_), .Y(_1772_) );
NAND3X1 NAND3X1_354 ( .gnd(gnd), .vdd(vdd), .A(_1580_), .B(_1772_), .C(_1766_), .Y(_1773_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1765_), .B(_1762_), .C(_1767_), .Y(_1774_) );
NAND3X1 NAND3X1_355 ( .gnd(gnd), .vdd(vdd), .A(_1734_), .B(_1770_), .C(_1771_), .Y(_1775_) );
NAND3X1 NAND3X1_356 ( .gnd(gnd), .vdd(vdd), .A(_1585_), .B(_1775_), .C(_1774_), .Y(_1776_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1776_), .B(_1773_), .Y(_1777_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(_3715_), .Y(_1778_) );
XNOR2X1 XNOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1778_), .B(bloque_datos[39]), .Y(_1779_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_1779_), .Y(_1780_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_1779_), .B(_1049_), .Y(_1781_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1781_), .B(_1780_), .C(_1777_), .Y(_1782_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_1773_), .B(_1776_), .Y(_1783_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_1779_), .B(_1049_), .Y(_1784_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_1779_), .Y(_1785_) );
NAND3X1 NAND3X1_357 ( .gnd(gnd), .vdd(vdd), .A(_1784_), .B(_1785_), .C(_1783_), .Y(_1786_) );
NAND3X1 NAND3X1_358 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .B(_1782_), .C(_1786_), .Y(_1787_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .B(_1061_), .C(_1054_), .Y(_1788_) );
AOI21X1 AOI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1784_), .B(_1785_), .C(_1783_), .Y(_1789_) );
NOR3X1 NOR3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1780_), .B(_1781_), .C(_1777_), .Y(_1790_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .B(_1790_), .C(_1788_), .Y(_1791_) );
NAND3X1 NAND3X1_359 ( .gnd(gnd), .vdd(vdd), .A(_1595_), .B(_1787_), .C(_1791_), .Y(_1792_) );
NAND3X1 NAND3X1_360 ( .gnd(gnd), .vdd(vdd), .A(_1788_), .B(_1782_), .C(_1786_), .Y(_1793_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .B(_1790_), .C(_1733_), .Y(_1794_) );
NAND3X1 NAND3X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1597_), .B(_1793_), .C(_1794_), .Y(_1795_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(_1795_), .Y(_1796_) );
XNOR2X1 XNOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_3725_), .B(bloque_datos[55]), .Y(_1797_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .B(_1084_), .Y(_1798_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_1797_), .Y(_1799_) );
AOI21X1 AOI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1799_), .B(_1798_), .C(_1796_), .Y(_1800_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(_1795_), .Y(_1801_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_1797_), .Y(_1802_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .B(_1084_), .Y(_1803_) );
NOR3X1 NOR3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(_1802_), .C(_1801_), .Y(_1804_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1800_), .B(_1804_), .C(_1732_), .Y(_1805_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1094_), .B(_1096_), .C(_1089_), .Y(_1806_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(_1802_), .C(_1801_), .Y(_1807_) );
NAND3X1 NAND3X1_362 ( .gnd(gnd), .vdd(vdd), .A(_1799_), .B(_1798_), .C(_1796_), .Y(_1808_) );
NAND3X1 NAND3X1_363 ( .gnd(gnd), .vdd(vdd), .A(_1807_), .B(_1806_), .C(_1808_), .Y(_1809_) );
NAND3X1 NAND3X1_364 ( .gnd(gnd), .vdd(vdd), .A(_1731_), .B(_1809_), .C(_1805_), .Y(_1810_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1800_), .B(_1804_), .C(_1806_), .Y(_1811_) );
NAND3X1 NAND3X1_365 ( .gnd(gnd), .vdd(vdd), .A(_1732_), .B(_1807_), .C(_1808_), .Y(_1812_) );
NAND3X1 NAND3X1_366 ( .gnd(gnd), .vdd(vdd), .A(_1730_), .B(_1812_), .C(_1811_), .Y(_1813_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .B(_1813_), .Y(_1814_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_3731_), .B(_3737_), .C(bloque_datos_71_bF_buf3_), .Y(_1815_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf2_), .Y(_1816_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_3733_), .B(_3736_), .C(_3732_), .Y(_1817_) );
NAND3X1 NAND3X1_367 ( .gnd(gnd), .vdd(vdd), .A(_3662_), .B(_3730_), .C(_3727_), .Y(_1818_) );
NAND3X1 NAND3X1_368 ( .gnd(gnd), .vdd(vdd), .A(_1816_), .B(_1817_), .C(_1818_), .Y(_1819_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1819_), .B(_1815_), .Y(_1820_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_1820_), .B(_1122_), .Y(_1821_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .B(_1820_), .Y(_1822_) );
AOI21X1 AOI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1821_), .B(_1822_), .C(_1814_), .Y(_1823_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .B(_1813_), .Y(_1824_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .B(_1820_), .Y(_1825_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_1820_), .B(_1122_), .Y(_1826_) );
NOR3X1 NOR3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1826_), .B(_1825_), .C(_1824_), .Y(_1827_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1823_), .B(_1827_), .C(_1729_), .Y(_1828_) );
AOI21X1 AOI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_970_), .C(_1133_), .Y(_1829_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1826_), .B(_1825_), .C(_1824_), .Y(_1830_) );
NAND3X1 NAND3X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1821_), .B(_1822_), .C(_1814_), .Y(_1831_) );
NAND3X1 NAND3X1_370 ( .gnd(gnd), .vdd(vdd), .A(_1829_), .B(_1830_), .C(_1831_), .Y(_1832_) );
AOI21X1 AOI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1832_), .B(_1828_), .C(_1728_), .Y(_1833_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(_1728_), .Y(_1834_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1823_), .B(_1827_), .C(_1829_), .Y(_1835_) );
NAND3X1 NAND3X1_371 ( .gnd(gnd), .vdd(vdd), .A(_1830_), .B(_1729_), .C(_1831_), .Y(_1836_) );
AOI21X1 AOI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1836_), .B(_1835_), .C(_1834_), .Y(_1837_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_1833_), .B(_1837_), .Y(_1838_) );
NAND3X1 NAND3X1_372 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf3_), .B(_3747_), .C(_3751_), .Y(_1839_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf2_), .Y(_1840_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .B(_3746_), .C(_1840_), .Y(_1841_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_1841_), .Y(_1842_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(_1164_), .Y(_1843_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1164_), .B(_1842_), .Y(_1844_) );
NAND3X1 NAND3X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1843_), .B(_1844_), .C(_1838_), .Y(_1845_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1833_), .B(_1837_), .Y(_1846_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1164_), .B(_1842_), .Y(_1847_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(_1164_), .Y(_1848_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_1847_), .C(_1846_), .Y(_1849_) );
NAND3X1 NAND3X1_374 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(_1727_), .C(_1845_), .Y(_1850_) );
AOI21X1 AOI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1172_), .B(_968_), .C(_1175_), .Y(_1851_) );
NOR3X1 NOR3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_1847_), .C(_1846_), .Y(_1852_) );
AOI21X1 AOI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1844_), .B(_1843_), .C(_1838_), .Y(_1853_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1852_), .B(_1853_), .C(_1851_), .Y(_1854_) );
AOI21X1 AOI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1850_), .B(_1854_), .C(_1726_), .Y(_1855_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(_1726_), .Y(_1856_) );
NAND3X1 NAND3X1_375 ( .gnd(gnd), .vdd(vdd), .A(_1851_), .B(_1849_), .C(_1845_), .Y(_1857_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1852_), .B(_1853_), .C(_1727_), .Y(_1858_) );
AOI21X1 AOI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1857_), .B(_1858_), .C(_1856_), .Y(_1859_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(_1859_), .Y(_1860_) );
NAND3X1 NAND3X1_376 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_135_), .B(_3759_), .C(_3762_), .Y(_1861_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_135_), .Y(_1862_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_3760_), .B(_3758_), .C(_1862_), .Y(_1863_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_1861_), .B(_1863_), .Y(_1864_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1864_), .B(_1205_), .Y(_1865_) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1864_), .B(_1205_), .Y(_1866_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_1866_), .Y(_1867_) );
NOR3X1 NOR3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .B(_1865_), .C(_1860_), .Y(_1868_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(_1859_), .Y(_1869_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(_1865_), .Y(_1870_) );
AOI21X1 AOI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1866_), .B(_1870_), .C(_1869_), .Y(_1871_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1868_), .B(_1871_), .C(_1725_), .Y(_1872_) );
NAND3X1 NAND3X1_377 ( .gnd(gnd), .vdd(vdd), .A(_1866_), .B(_1870_), .C(_1869_), .Y(_1873_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .B(_1865_), .C(_1860_), .Y(_1874_) );
NAND3X1 NAND3X1_378 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_1874_), .C(_1873_), .Y(_1875_) );
AOI21X1 AOI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1875_), .B(_1872_), .C(_1639_), .Y(_1876_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .Y(_1877_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1868_), .B(_1871_), .C(_1724_), .Y(_1878_) );
NAND3X1 NAND3X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1874_), .B(_1873_), .C(_1725_), .Y(_1879_) );
AOI21X1 AOI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1879_), .B(_1878_), .C(_1877_), .Y(_1880_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1876_), .B(_1880_), .C(_1723_), .Y(_1881_) );
NAND3X1 NAND3X1_380 ( .gnd(gnd), .vdd(vdd), .A(_1877_), .B(_1879_), .C(_1878_), .Y(_1882_) );
NAND3X1 NAND3X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(_1875_), .C(_1872_), .Y(_1883_) );
NAND3X1 NAND3X1_382 ( .gnd(gnd), .vdd(vdd), .A(_1245_), .B(_1882_), .C(_1883_), .Y(_1884_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1884_), .B(_1881_), .Y(_1885_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_1278_), .C(_1885_), .Y(_1886_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(_3771_), .Y(_1887_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1255_), .B(_1257_), .C(_1250_), .Y(_1888_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(_1888_), .Y(_1889_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_1881_), .B(_1884_), .Y(_1890_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_3768_), .B(_1887_), .C(_1890_), .D(_1889_), .Y(_1891_) );
NAND3X1 NAND3X1_383 ( .gnd(gnd), .vdd(vdd), .A(_1648_), .B(_1886_), .C(_1891_), .Y(_1892_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(_1648_), .Y(_1893_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1889_), .B(_1890_), .Y(_1894_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_3768_), .B(_1887_), .Y(_1895_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1885_), .B(_1888_), .C(_1895_), .Y(_1896_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1894_), .B(_1896_), .C(_1893_), .Y(_1897_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_1892_), .B(_1897_), .Y(_1898_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_151_), .Y(_1899_) );
AOI21X1 AOI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_150_), .B(_1281_), .C(_1899_), .Y(_1900_) );
NOR3X1 NOR3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(module_0_W_151_), .C(_1286_), .Y(_1901_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1900_), .B(_1901_), .C(_1898_), .Y(_1902_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1897_), .B(_1892_), .Y(_1903_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1283_), .C(module_0_W_151_), .Y(_1904_) );
NAND3X1 NAND3X1_384 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_150_), .B(_1899_), .C(_1281_), .Y(_1905_) );
NAND3X1 NAND3X1_385 ( .gnd(gnd), .vdd(vdd), .A(_1904_), .B(_1905_), .C(_1903_), .Y(_1906_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .B(_1906_), .Y(_1907_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(_1292_), .C(_1907_), .Y(_1908_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_960_), .B(_1313_), .C(_1295_), .Y(_1909_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(_1909_), .Y(_1910_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1906_), .B(_1902_), .Y(_1911_) );
AOI21X1 AOI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1911_), .B(_1910_), .C(_3783_), .Y(_1912_) );
NAND3X1 NAND3X1_386 ( .gnd(gnd), .vdd(vdd), .A(_1722_), .B(_1908_), .C(_1912_), .Y(_1913_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1911_), .B(_1910_), .Y(_1914_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(_3783_), .Y(_1915_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1907_), .B(_1909_), .C(_1915_), .Y(_1916_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(_1914_), .C(_1661_), .Y(_1917_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1913_), .B(_1917_), .Y(_1918_) );
AOI21X1 AOI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1719_), .B(_1721_), .C(_1918_), .Y(_1919_) );
NAND3X1 NAND3X1_387 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_166_), .B(module_0_W_167_), .C(_1316_), .Y(_1920_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1321_), .B(_1318_), .C(_1720_), .Y(_1921_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1913_), .B(_1917_), .C(_1921_), .D(_1920_), .Y(_1922_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1922_), .B(_1919_), .Y(_1923_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1347_), .B(_1327_), .C(_1923_), .Y(_1924_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_958_), .C(_1330_), .Y(_1925_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(_1925_), .Y(_1926_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1920_), .B(_1921_), .Y(_1927_) );
XNOR2X1 XNOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1927_), .B(_1918_), .Y(_1928_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_3791_), .B(_3793_), .C(_1928_), .D(_1926_), .Y(_1929_) );
NAND3X1 NAND3X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1718_), .B(_1924_), .C(_1929_), .Y(_1930_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .B(_1926_), .Y(_1931_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1923_), .B(_1925_), .C(_3794_), .Y(_1932_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1931_), .B(_1932_), .C(_1671_), .Y(_1933_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_1933_), .Y(_1934_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_183_), .Y(_1935_) );
AOI21X1 AOI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_182_), .B(_1351_), .C(_1935_), .Y(_1936_) );
NOR3X1 NOR3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1353_), .B(module_0_W_183_), .C(_1356_), .Y(_1937_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1936_), .B(_1937_), .C(_1934_), .Y(_1938_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1933_), .B(_1930_), .Y(_1939_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .B(_1353_), .C(module_0_W_183_), .Y(_1940_) );
NAND3X1 NAND3X1_389 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_182_), .B(_1935_), .C(_1351_), .Y(_1941_) );
NAND3X1 NAND3X1_390 ( .gnd(gnd), .vdd(vdd), .A(_1940_), .B(_1941_), .C(_1939_), .Y(_1942_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1942_), .B(_1938_), .Y(_1943_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1943_), .B(_1717_), .Y(_1944_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(_1942_), .Y(_1945_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1945_), .B(_1716_), .C(_376_), .Y(_1946_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_1944_), .C(module_0_W_199_), .Y(_1947_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_199_), .Y(_1948_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .B(_1385_), .C(_1945_), .Y(_1950_) );
AOI21X1 AOI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1943_), .B(_1717_), .C(_3808_), .Y(_1951_) );
NAND3X1 NAND3X1_391 ( .gnd(gnd), .vdd(vdd), .A(_1948_), .B(_1950_), .C(_1951_), .Y(_1952_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1952_), .B(_1947_), .Y(_1953_) );
NOR3X1 NOR3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1385_), .B(_1387_), .C(_1386_), .Y(_1954_) );
NOR3X1 NOR3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_1392_), .C(_1954_), .Y(_1955_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1955_), .B(_1391_), .C(_1680_), .Y(_1956_) );
INVX2 INVX2_62 ( .gnd(gnd), .vdd(vdd), .A(_1680_), .Y(_1957_) );
NAND3X1 NAND3X1_392 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_198_), .B(_1957_), .C(_1389_), .Y(_1958_) );
NAND3X1 NAND3X1_393 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .B(_1958_), .C(_1953_), .Y(_1959_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_1947_), .B(_1952_), .Y(_1961_) );
AOI21X1 AOI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_198_), .B(_1389_), .C(_1957_), .Y(_1962_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(_1958_), .Y(_1963_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1963_), .B(_1962_), .C(_1961_), .Y(_1964_) );
AOI21X1 AOI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1959_), .B(_1964_), .C(_1715_), .Y(_1965_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(_951_), .C(_1402_), .Y(_1966_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1959_), .B(_1964_), .Y(_1967_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1967_), .B(_1966_), .C(_3823_), .Y(_1968_) );
NOR3X1 NOR3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1965_), .B(_1691_), .C(_1968_), .Y(_1969_) );
INVX2 INVX2_63 ( .gnd(gnd), .vdd(vdd), .A(_1691_), .Y(_1970_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(_1965_), .Y(_1972_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_1964_), .B(_1959_), .Y(_1973_) );
AOI21X1 AOI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1715_), .B(_1973_), .C(_3826_), .Y(_1974_) );
AOI21X1 AOI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1972_), .B(_1974_), .C(_1970_), .Y(_1975_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1969_), .B(_1975_), .Y(_1976_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_215_), .Y(_1977_) );
AOI21X1 AOI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_214_), .B(_1425_), .C(_1977_), .Y(_1978_) );
NOR3X1 NOR3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1427_), .B(module_0_W_215_), .C(_1430_), .Y(_1979_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1978_), .B(_1979_), .C(_1976_), .Y(_1980_) );
NAND3X1 NAND3X1_394 ( .gnd(gnd), .vdd(vdd), .A(_1970_), .B(_1972_), .C(_1974_), .Y(_1981_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1968_), .B(_1965_), .C(_1691_), .Y(_1983_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1983_), .B(_1981_), .Y(_1984_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1430_), .B(_1427_), .C(module_0_W_215_), .Y(_1985_) );
NAND3X1 NAND3X1_395 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_214_), .B(_1977_), .C(_1425_), .Y(_1986_) );
NAND3X1 NAND3X1_396 ( .gnd(gnd), .vdd(vdd), .A(_1985_), .B(_1986_), .C(_1984_), .Y(_1987_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_1980_), .B(_1987_), .Y(_1988_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_1458_), .B(_1436_), .C(_1988_), .Y(_1989_) );
AOI21X1 AOI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1440_), .B(_1438_), .C(_1458_), .Y(_1990_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1987_), .B(_1980_), .Y(_1991_) );
AOI21X1 AOI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_1991_), .C(_3835_), .Y(_1992_) );
NAND3X1 NAND3X1_397 ( .gnd(gnd), .vdd(vdd), .A(_1714_), .B(_1992_), .C(_1989_), .Y(_1994_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_1991_), .Y(_1995_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(_3835_), .Y(_1996_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_1459_), .B(_948_), .C(_1439_), .Y(_1997_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_1988_), .B(_1997_), .C(_1996_), .Y(_1998_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_1998_), .B(_1995_), .C(_1701_), .Y(_1999_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_1999_), .B(_1994_), .Y(_2000_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_231_), .Y(_2001_) );
AOI21X1 AOI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_230_), .B(_1462_), .C(_2001_), .Y(_2002_) );
NOR3X1 NOR3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(module_0_W_231_), .C(_1467_), .Y(_2003_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_2002_), .B(_2003_), .C(_2000_), .Y(_2005_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1994_), .B(_1999_), .Y(_2006_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1467_), .B(_1464_), .C(module_0_W_231_), .Y(_2007_) );
NAND3X1 NAND3X1_398 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_230_), .B(_2001_), .C(_1462_), .Y(_2008_) );
NAND3X1 NAND3X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2007_), .B(_2008_), .C(_2006_), .Y(_2009_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .B(_2009_), .Y(_2010_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1495_), .B(_1473_), .C(_2010_), .Y(_2011_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1496_), .B(_942_), .C(_1476_), .Y(_2012_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .Y(_2013_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_2009_), .B(_2005_), .Y(_2014_) );
AOI21X1 AOI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_2014_), .B(_2013_), .C(_3848_), .Y(_2016_) );
NAND3X1 NAND3X1_400 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_247_), .B(_2011_), .C(_2016_), .Y(_2017_) );
INVX2 INVX2_64 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_247_), .Y(_2018_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_2014_), .B(_2013_), .Y(_2019_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(_3848_), .Y(_2020_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_2010_), .B(_2012_), .C(_2020_), .Y(_2021_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_2021_), .B(_2019_), .C(_2018_), .Y(_2022_) );
NAND3X1 NAND3X1_401 ( .gnd(gnd), .vdd(vdd), .A(_2017_), .B(_2022_), .C(_1500_), .Y(_2023_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1501_), .B(_1504_), .Y(_2024_) );
NOR3X1 NOR3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_2019_), .B(_2018_), .C(_2021_), .Y(_2025_) );
AOI21X1 AOI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_2011_), .B(_2016_), .C(module_0_W_247_), .Y(_2027_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .B(_2027_), .C(_2024_), .Y(_2028_) );
NAND3X1 NAND3X1_402 ( .gnd(gnd), .vdd(vdd), .A(_1713_), .B(_2023_), .C(_2028_), .Y(_2029_) );
NAND3X1 NAND3X1_403 ( .gnd(gnd), .vdd(vdd), .A(_2018_), .B(_2011_), .C(_2016_), .Y(_2030_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_2021_), .B(_2019_), .C(module_0_W_247_), .Y(_2031_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_246_), .B(_1499_), .C(_2031_), .D(_2030_), .Y(_2032_) );
AOI21X1 AOI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_2017_), .B(_2022_), .C(_1500_), .Y(_2033_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2033_), .B(_2032_), .C(_1712_), .Y(_2034_) );
NAND3X1 NAND3X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2029_), .B(_2034_), .C(_1537_), .Y(_2035_) );
AOI21X1 AOI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1500_), .B(_1505_), .C(_917_), .Y(_2036_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_2036_), .B(_940_), .C(_1512_), .Y(_2038_) );
NOR3X1 NOR3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_2032_), .B(_1712_), .C(_2033_), .Y(_2039_) );
AOI21X1 AOI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_2023_), .B(_2028_), .C(_1713_), .Y(_2040_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_2039_), .B(_2040_), .C(_2038_), .Y(_2041_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_2041_), .B(_2035_), .Y(_2042_) );
NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_2042_), .B(_1535_), .Y(_2043_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_2039_), .B(_2040_), .C(_1537_), .Y(_2044_) );
NAND3X1 NAND3X1_405 ( .gnd(gnd), .vdd(vdd), .A(_2029_), .B(_2034_), .C(_2038_), .Y(_2045_) );
NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_2045_), .B(_2044_), .Y(_2046_) );
NAND3X1 NAND3X1_406 ( .gnd(gnd), .vdd(vdd), .A(_939_), .B(_2046_), .C(_1532_), .Y(_2047_) );
NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_2047_), .B(_2043_), .Y(module_0_H_7_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_248_), .B(_464_), .Y(_2049_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(_2049_), .Y(_2050_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_458_), .C(module_0_W_248_), .Y(_2051_) );
NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_2051_), .B(_2050_), .Y(module_0_H_16_) );
XNOR2X1 XNOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(module_0_W_249_), .Y(_2052_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(_2052_), .Y(_2053_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_248_), .B(_464_), .C(_2053_), .Y(_2054_) );
INVX2 INVX2_65 ( .gnd(gnd), .vdd(vdd), .A(_2054_), .Y(_2055_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_2050_), .B(_2053_), .Y(_2056_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_2056_), .B(_2055_), .Y(module_0_H_17_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_249_), .B(_934_), .Y(_2058_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(_2058_), .Y(_2059_) );
NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_250_), .B(_1526_), .Y(_2060_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_1526_), .B(module_0_W_250_), .Y(_2061_) );
AOI21X1 AOI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(_2061_), .C(_2059_), .Y(_2062_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(_2062_), .Y(_2063_) );
NAND3X1 NAND3X1_407 ( .gnd(gnd), .vdd(vdd), .A(_2059_), .B(_2060_), .C(_2061_), .Y(_2064_) );
NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_2064_), .B(_2063_), .Y(_2065_) );
XNOR2X1 XNOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .B(_2055_), .Y(module_0_H_18_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2062_), .B(_2054_), .C(_2064_), .Y(_2067_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_250_), .B(_1527_), .Y(_2068_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_251_), .Y(_2069_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(_1708_), .C(_2069_), .Y(_2070_) );
NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_251_), .B(_1712_), .Y(_2071_) );
NAND3X1 NAND3X1_408 ( .gnd(gnd), .vdd(vdd), .A(_2068_), .B(_2070_), .C(_2071_), .Y(_2072_) );
AOI21X1 AOI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_2070_), .B(_2071_), .C(_2068_), .Y(_2073_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(_2073_), .Y(_2074_) );
NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_2072_), .B(_2074_), .Y(_2075_) );
XNOR2X1 XNOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_2075_), .B(_2067_), .Y(module_0_H_19_) );
AOI21X1 AOI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_2067_), .B(_2072_), .C(_2073_), .Y(_2077_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1706_), .C(_1704_), .Y(_2078_) );
INVX2 INVX2_66 ( .gnd(gnd), .vdd(vdd), .A(_1703_), .Y(_2079_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1693_), .B(_1692_), .C(_1483_), .Y(_2080_) );
AOI21X1 AOI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_2080_), .B(_1539_), .C(_1694_), .Y(_2081_) );
NOR3X1 NOR3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1446_), .B(_1682_), .C(_1685_), .Y(_2082_) );
AOI21X1 AOI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1686_), .B(_1689_), .C(_2082_), .Y(_2083_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1678_), .B(_1675_), .C(_1673_), .Y(_2084_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(_1672_), .Y(_2085_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_1663_), .B(_1546_), .Y(_2086_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .B(_1544_), .C(_2086_), .Y(_2088_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1547_), .B(_1722_), .Y(_2089_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1650_), .B(_1651_), .C(_1336_), .Y(_2090_) );
AOI21X1 AOI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_2090_), .B(_1548_), .C(_1652_), .Y(_2091_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1646_), .B(_1550_), .C(_1642_), .Y(_2092_) );
INVX2 INVX2_67 ( .gnd(gnd), .vdd(vdd), .A(_2092_), .Y(_2093_) );
NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_139_), .B(_1639_), .Y(_2094_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(_1632_), .Y(_2095_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .Y(_2096_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf3_), .Y(_2097_) );
XNOR2X1 XNOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_2592_), .Y(_2099_) );
NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(_1626_), .Y(_2100_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_2120_), .Y(_2101_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(_1555_), .Y(_2102_) );
AOI21X1 AOI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .B(_1607_), .C(_1183_), .Y(_2103_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_2102_), .B(_2103_), .C(_1610_), .Y(_2104_) );
XNOR2X1 XNOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_2087_), .Y(_2105_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_1146_), .B(_513_), .C(_1149_), .Y(_2106_) );
AOI21X1 AOI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1600_), .B(_2106_), .C(_1599_), .Y(_2107_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(_1596_), .Y(_2108_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf4_), .Y(_2110_) );
AOI21X1 AOI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1593_), .B(_1591_), .C(_1588_), .Y(_2111_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf2_), .B(_1585_), .Y(_2112_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf4_), .Y(_2113_) );
XNOR2X1 XNOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_3978_), .B(_2026_), .Y(_2114_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(_2114_), .Y(_2115_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_1579_), .B(_1561_), .C(_1577_), .Y(_2116_) );
XNOR2X1 XNOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_3954_), .B(_2004_), .Y(_2117_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(_2117_), .Y(_2118_) );
AOI21X1 AOI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1033_), .B(_491_), .C(_1037_), .Y(_2119_) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_2119_), .B(_1571_), .C(_1569_), .Y(_2121_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_28_), .Y(_2122_) );
XNOR2X1 XNOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_0_), .B(module_0_W_12_), .Y(_2123_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_2123_), .B(module_0_W_8_), .Y(_2124_) );
NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_2122_), .B(_2124_), .Y(_2125_) );
XNOR2X1 XNOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_2123_), .B(module_0_W_8_), .Y(_2126_) );
NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_28_), .B(_2126_), .Y(_2127_) );
NAND3X1 NAND3X1_409 ( .gnd(gnd), .vdd(vdd), .A(_1565_), .B(_2127_), .C(_2125_), .Y(_2128_) );
AOI21X1 AOI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_2127_), .B(_2125_), .C(_1565_), .Y(_2129_) );
INVX2 INVX2_68 ( .gnd(gnd), .vdd(vdd), .A(_2129_), .Y(_2130_) );
AOI21X1 AOI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_2128_), .B(_2130_), .C(_2121_), .Y(_2132_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .Y(_2133_) );
AOI21X1 AOI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1570_), .B(_1564_), .C(_2133_), .Y(_2134_) );
INVX2 INVX2_69 ( .gnd(gnd), .vdd(vdd), .A(_2128_), .Y(_2135_) );
NOR3X1 NOR3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_2134_), .B(_2129_), .C(_2135_), .Y(_2136_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2136_), .B(_2132_), .C(_2118_), .Y(_2137_) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_2135_), .B(_2129_), .C(_2134_), .Y(_2138_) );
NAND3X1 NAND3X1_410 ( .gnd(gnd), .vdd(vdd), .A(_2121_), .B(_2128_), .C(_2130_), .Y(_2139_) );
NAND3X1 NAND3X1_411 ( .gnd(gnd), .vdd(vdd), .A(_2117_), .B(_2139_), .C(_2138_), .Y(_2140_) );
NAND3X1 NAND3X1_412 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf3_), .B(_2140_), .C(_2137_), .Y(_2141_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf2_), .Y(_2143_) );
NAND3X1 NAND3X1_413 ( .gnd(gnd), .vdd(vdd), .A(_2118_), .B(_2139_), .C(_2138_), .Y(_2144_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_2136_), .B(_2132_), .C(_2117_), .Y(_2145_) );
NAND3X1 NAND3X1_414 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(_2144_), .C(_2145_), .Y(_2146_) );
NAND3X1 NAND3X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1573_), .B(_2141_), .C(_2146_), .Y(_2147_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(_1573_), .Y(_2148_) );
NAND3X1 NAND3X1_416 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(_2140_), .C(_2137_), .Y(_2149_) );
NAND3X1 NAND3X1_417 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf1_), .B(_2144_), .C(_2145_), .Y(_2150_) );
NAND3X1 NAND3X1_418 ( .gnd(gnd), .vdd(vdd), .A(_2148_), .B(_2149_), .C(_2150_), .Y(_2151_) );
AOI21X1 AOI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_2147_), .B(_2151_), .C(_2116_), .Y(_2152_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(_1577_), .Y(_2154_) );
AOI21X1 AOI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1578_), .B(_1584_), .C(_2154_), .Y(_2155_) );
AOI21X1 AOI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_2149_), .B(_2150_), .C(_2148_), .Y(_2156_) );
AOI21X1 AOI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_2141_), .B(_2146_), .C(_1573_), .Y(_2157_) );
NOR3X1 NOR3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_2156_), .B(_2155_), .C(_2157_), .Y(_2158_) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_2158_), .B(_2152_), .C(_2115_), .Y(_2159_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_2156_), .B(_2157_), .C(_2155_), .Y(_2160_) );
NAND3X1 NAND3X1_419 ( .gnd(gnd), .vdd(vdd), .A(_2147_), .B(_2151_), .C(_2116_), .Y(_2161_) );
NAND3X1 NAND3X1_420 ( .gnd(gnd), .vdd(vdd), .A(_2114_), .B(_2160_), .C(_2161_), .Y(_2162_) );
NAND3X1 NAND3X1_421 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(_2162_), .C(_2159_), .Y(_2163_) );
NAND3X1 NAND3X1_422 ( .gnd(gnd), .vdd(vdd), .A(_2115_), .B(_2160_), .C(_2161_), .Y(_2165_) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_2158_), .B(_2152_), .C(_2114_), .Y(_2166_) );
NAND3X1 NAND3X1_423 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf3_), .B(_2165_), .C(_2166_), .Y(_2167_) );
AOI21X1 AOI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(_2167_), .C(_2112_), .Y(_2168_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(_2112_), .Y(_2169_) );
NAND3X1 NAND3X1_424 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf2_), .B(_2162_), .C(_2159_), .Y(_2170_) );
NAND3X1 NAND3X1_425 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(_2165_), .C(_2166_), .Y(_2171_) );
AOI21X1 AOI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_2170_), .B(_2171_), .C(_2169_), .Y(_2172_) );
OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_2168_), .B(_2172_), .C(_2111_), .Y(_2173_) );
OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_1559_), .B(_1589_), .C(_1592_), .Y(_2174_) );
NAND3X1 NAND3X1_426 ( .gnd(gnd), .vdd(vdd), .A(_2169_), .B(_2170_), .C(_2171_), .Y(_2176_) );
NAND3X1 NAND3X1_427 ( .gnd(gnd), .vdd(vdd), .A(_2112_), .B(_2163_), .C(_2167_), .Y(_2177_) );
NAND3X1 NAND3X1_428 ( .gnd(gnd), .vdd(vdd), .A(_2176_), .B(_2177_), .C(_2174_), .Y(_2178_) );
XNOR2X1 XNOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_2057_), .Y(_2179_) );
NAND3X1 NAND3X1_429 ( .gnd(gnd), .vdd(vdd), .A(_2179_), .B(_2178_), .C(_2173_), .Y(_2180_) );
AOI21X1 AOI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_2176_), .B(_2177_), .C(_2174_), .Y(_2181_) );
NOR3X1 NOR3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_2168_), .B(_2172_), .C(_2111_), .Y(_2182_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(_2179_), .Y(_2183_) );
OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_2182_), .B(_2181_), .C(_2183_), .Y(_2184_) );
NAND3X1 NAND3X1_430 ( .gnd(gnd), .vdd(vdd), .A(_2110_), .B(_2180_), .C(_2184_), .Y(_2185_) );
NAND3X1 NAND3X1_431 ( .gnd(gnd), .vdd(vdd), .A(_2183_), .B(_2178_), .C(_2173_), .Y(_2187_) );
OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_2182_), .B(_2181_), .C(_2179_), .Y(_2188_) );
NAND3X1 NAND3X1_432 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf3_), .B(_2187_), .C(_2188_), .Y(_2189_) );
AOI21X1 AOI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_2185_), .B(_2189_), .C(_2108_), .Y(_2190_) );
NAND3X1 NAND3X1_433 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf2_), .B(_2180_), .C(_2184_), .Y(_2191_) );
NAND3X1 NAND3X1_434 ( .gnd(gnd), .vdd(vdd), .A(_2110_), .B(_2187_), .C(_2188_), .Y(_2192_) );
AOI21X1 AOI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_2191_), .B(_2192_), .C(_1596_), .Y(_2193_) );
OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_2190_), .B(_2193_), .C(_2107_), .Y(_2194_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(_1599_), .Y(_2195_) );
OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_1556_), .B(_1601_), .C(_2195_), .Y(_2196_) );
NAND3X1 NAND3X1_435 ( .gnd(gnd), .vdd(vdd), .A(_1596_), .B(_2191_), .C(_2192_), .Y(_2198_) );
NAND3X1 NAND3X1_436 ( .gnd(gnd), .vdd(vdd), .A(_2108_), .B(_2185_), .C(_2189_), .Y(_2199_) );
NAND3X1 NAND3X1_437 ( .gnd(gnd), .vdd(vdd), .A(_2198_), .B(_2199_), .C(_2196_), .Y(_2200_) );
NAND3X1 NAND3X1_438 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .B(_2194_), .C(_2200_), .Y(_2201_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .Y(_2202_) );
AOI21X1 AOI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_2198_), .B(_2199_), .C(_2196_), .Y(_2203_) );
NOR3X1 NOR3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_2190_), .B(_2193_), .C(_2107_), .Y(_2204_) );
OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_2204_), .B(_2203_), .C(_2202_), .Y(_2205_) );
NAND3X1 NAND3X1_439 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf3_), .B(_2201_), .C(_2205_), .Y(_2206_) );
INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf2_), .Y(_2207_) );
NAND3X1 NAND3X1_440 ( .gnd(gnd), .vdd(vdd), .A(_2202_), .B(_2194_), .C(_2200_), .Y(_2209_) );
OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2204_), .B(_2203_), .C(_2105_), .Y(_2210_) );
NAND3X1 NAND3X1_441 ( .gnd(gnd), .vdd(vdd), .A(_2207_), .B(_2209_), .C(_2210_), .Y(_2211_) );
NAND3X1 NAND3X1_442 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(_2206_), .C(_2211_), .Y(_2212_) );
INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .Y(_2213_) );
NAND3X1 NAND3X1_443 ( .gnd(gnd), .vdd(vdd), .A(_2207_), .B(_2201_), .C(_2205_), .Y(_2214_) );
NAND3X1 NAND3X1_444 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf1_), .B(_2209_), .C(_2210_), .Y(_2215_) );
NAND3X1 NAND3X1_445 ( .gnd(gnd), .vdd(vdd), .A(_2213_), .B(_2214_), .C(_2215_), .Y(_2216_) );
AOI21X1 AOI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_2212_), .B(_2216_), .C(_2104_), .Y(_2217_) );
AOI21X1 AOI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_1612_), .B(_1611_), .C(_1186_), .Y(_2218_) );
AOI21X1 AOI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_1555_), .B(_1613_), .C(_2218_), .Y(_2220_) );
AOI21X1 AOI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_2214_), .B(_2215_), .C(_2213_), .Y(_2221_) );
AOI21X1 AOI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_2206_), .B(_2211_), .C(_1611_), .Y(_2222_) );
NOR3X1 NOR3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_2221_), .B(_2222_), .C(_2220_), .Y(_2223_) );
OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_2223_), .B(_2217_), .C(_2101_), .Y(_2224_) );
INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .Y(_2225_) );
OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_2221_), .B(_2222_), .C(_2220_), .Y(_2226_) );
NAND3X1 NAND3X1_446 ( .gnd(gnd), .vdd(vdd), .A(_2212_), .B(_2216_), .C(_2104_), .Y(_2227_) );
NAND3X1 NAND3X1_447 ( .gnd(gnd), .vdd(vdd), .A(_2225_), .B(_2226_), .C(_2227_), .Y(_2228_) );
NAND3X1 NAND3X1_448 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf4_), .B(_2228_), .C(_2224_), .Y(_2229_) );
INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf3_), .Y(_2231_) );
NAND3X1 NAND3X1_449 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .B(_2226_), .C(_2227_), .Y(_2232_) );
OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_2223_), .B(_2217_), .C(_2225_), .Y(_2233_) );
NAND3X1 NAND3X1_450 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .B(_2232_), .C(_2233_), .Y(_2234_) );
NAND3X1 NAND3X1_451 ( .gnd(gnd), .vdd(vdd), .A(_1622_), .B(_2229_), .C(_2234_), .Y(_2235_) );
INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(_1622_), .Y(_2236_) );
NAND3X1 NAND3X1_452 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .B(_2228_), .C(_2224_), .Y(_2237_) );
NAND3X1 NAND3X1_453 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf2_), .B(_2232_), .C(_2233_), .Y(_2238_) );
NAND3X1 NAND3X1_454 ( .gnd(gnd), .vdd(vdd), .A(_2236_), .B(_2237_), .C(_2238_), .Y(_2239_) );
AOI21X1 AOI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_2235_), .B(_2239_), .C(_2100_), .Y(_2240_) );
INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .Y(_2242_) );
AOI21X1 AOI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1624_), .B(_1553_), .C(_2242_), .Y(_2243_) );
AOI21X1 AOI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_2237_), .B(_2238_), .C(_2236_), .Y(_2244_) );
AOI21X1 AOI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .B(_2234_), .C(_1622_), .Y(_2245_) );
NOR3X1 NOR3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_2244_), .B(_2243_), .C(_2245_), .Y(_2246_) );
OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_2246_), .B(_2240_), .C(_2099_), .Y(_2247_) );
INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(_2099_), .Y(_2248_) );
OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_2244_), .B(_2245_), .C(_2243_), .Y(_2249_) );
NAND3X1 NAND3X1_455 ( .gnd(gnd), .vdd(vdd), .A(_2235_), .B(_2239_), .C(_2100_), .Y(_2250_) );
NAND3X1 NAND3X1_456 ( .gnd(gnd), .vdd(vdd), .A(_2248_), .B(_2250_), .C(_2249_), .Y(_2251_) );
NAND3X1 NAND3X1_457 ( .gnd(gnd), .vdd(vdd), .A(_2097_), .B(_2251_), .C(_2247_), .Y(_2253_) );
NAND3X1 NAND3X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2099_), .B(_2250_), .C(_2249_), .Y(_2254_) );
OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_2246_), .B(_2240_), .C(_2248_), .Y(_2255_) );
NAND3X1 NAND3X1_459 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf2_), .B(_2254_), .C(_2255_), .Y(_2256_) );
AOI21X1 AOI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_2253_), .B(_2256_), .C(_2096_), .Y(_2257_) );
NAND3X1 NAND3X1_460 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf1_), .B(_2251_), .C(_2247_), .Y(_2258_) );
NAND3X1 NAND3X1_461 ( .gnd(gnd), .vdd(vdd), .A(_2097_), .B(_2254_), .C(_2255_), .Y(_2259_) );
AOI21X1 AOI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_2258_), .B(_2259_), .C(_1633_), .Y(_2260_) );
OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_2257_), .B(_2260_), .C(_2095_), .Y(_2261_) );
NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_1632_), .B(_1636_), .Y(_2262_) );
NAND3X1 NAND3X1_462 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .B(_2258_), .C(_2259_), .Y(_2264_) );
NAND3X1 NAND3X1_463 ( .gnd(gnd), .vdd(vdd), .A(_2096_), .B(_2253_), .C(_2256_), .Y(_2265_) );
NAND3X1 NAND3X1_464 ( .gnd(gnd), .vdd(vdd), .A(_2262_), .B(_2264_), .C(_2265_), .Y(_2266_) );
NAND3X1 NAND3X1_465 ( .gnd(gnd), .vdd(vdd), .A(_2570_), .B(_2266_), .C(_2261_), .Y(_2267_) );
AOI21X1 AOI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .B(_2265_), .C(_2262_), .Y(_2268_) );
NOR3X1 NOR3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_2260_), .B(_2095_), .C(_2257_), .Y(_2269_) );
OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_2269_), .B(_2268_), .C(_2186_), .Y(_2270_) );
NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2267_), .B(_2270_), .Y(_2271_) );
NAND3X1 NAND3X1_466 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_140_), .B(_292_), .C(_2271_), .Y(_2272_) );
INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_140_), .Y(_2273_) );
OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_2269_), .B(_2268_), .C(_2570_), .Y(_2275_) );
NAND3X1 NAND3X1_467 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(_2266_), .C(_2261_), .Y(_2276_) );
NAND3X1 NAND3X1_468 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(_2276_), .C(_2275_), .Y(_2277_) );
NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_2273_), .B(_2277_), .Y(_2278_) );
AOI21X1 AOI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2272_), .B(_2278_), .C(_2094_), .Y(_2279_) );
INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(_2094_), .Y(_2280_) );
NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_140_), .B(_2277_), .Y(_2281_) );
NAND3X1 NAND3X1_469 ( .gnd(gnd), .vdd(vdd), .A(_2273_), .B(_292_), .C(_2271_), .Y(_2282_) );
AOI21X1 AOI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_2281_), .B(_2282_), .C(_2280_), .Y(_2283_) );
OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2283_), .B(_2279_), .C(_2093_), .Y(_2284_) );
NAND3X1 NAND3X1_470 ( .gnd(gnd), .vdd(vdd), .A(_2280_), .B(_2281_), .C(_2282_), .Y(_2286_) );
NAND3X1 NAND3X1_471 ( .gnd(gnd), .vdd(vdd), .A(_2094_), .B(_2272_), .C(_2278_), .Y(_2287_) );
NAND3X1 NAND3X1_472 ( .gnd(gnd), .vdd(vdd), .A(_2092_), .B(_2286_), .C(_2287_), .Y(_2288_) );
NAND3X1 NAND3X1_473 ( .gnd(gnd), .vdd(vdd), .A(_2219_), .B(_2288_), .C(_2284_), .Y(_2289_) );
NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_2288_), .B(_2284_), .Y(_2290_) );
AOI21X1 AOI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_2537_), .B(_2290_), .C(_321_), .Y(_2291_) );
NAND3X1 NAND3X1_474 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_156_), .B(_2289_), .C(_2291_), .Y(_2292_) );
INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_156_), .Y(_2293_) );
AOI21X1 AOI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_2286_), .B(_2287_), .C(_2092_), .Y(_2294_) );
NOR3X1 NOR3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_2279_), .B(_2283_), .C(_2093_), .Y(_2295_) );
OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2295_), .B(_2294_), .C(_2537_), .Y(_2297_) );
NAND3X1 NAND3X1_475 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_2289_), .C(_2297_), .Y(_2298_) );
NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .B(_2298_), .Y(_2299_) );
AOI21X1 AOI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2292_), .B(_2299_), .C(_1653_), .Y(_2300_) );
NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_156_), .B(_2298_), .Y(_2301_) );
NAND3X1 NAND3X1_476 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .B(_2289_), .C(_2291_), .Y(_2302_) );
AOI21X1 AOI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_2302_), .B(_2301_), .C(_1651_), .Y(_2303_) );
OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2303_), .B(_2300_), .C(_2091_), .Y(_2304_) );
NAND3X1 NAND3X1_477 ( .gnd(gnd), .vdd(vdd), .A(_1335_), .B(_1649_), .C(_1653_), .Y(_2305_) );
OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .B(_1654_), .C(_2305_), .Y(_2306_) );
NAND3X1 NAND3X1_478 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .B(_2302_), .C(_2301_), .Y(_2308_) );
NAND3X1 NAND3X1_479 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_2292_), .C(_2299_), .Y(_2309_) );
NAND3X1 NAND3X1_480 ( .gnd(gnd), .vdd(vdd), .A(_2306_), .B(_2308_), .C(_2309_), .Y(_2310_) );
AOI21X1 AOI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2310_), .B(_2304_), .C(_2252_), .Y(_2311_) );
NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2310_), .B(_2304_), .Y(_2312_) );
OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_2312_), .B(_2504_), .C(_343_), .Y(_2313_) );
OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_2313_), .B(_2311_), .C(module_0_W_172_), .Y(_2314_) );
INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_172_), .Y(_2315_) );
NAND3X1 NAND3X1_481 ( .gnd(gnd), .vdd(vdd), .A(_2504_), .B(_2310_), .C(_2304_), .Y(_2316_) );
AOI21X1 AOI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_2308_), .B(_2309_), .C(_2306_), .Y(_2317_) );
NOR3X1 NOR3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_2300_), .B(_2091_), .C(_2303_), .Y(_2319_) );
OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_2319_), .B(_2317_), .C(_2252_), .Y(_2320_) );
NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_2316_), .B(_2320_), .Y(_2321_) );
NAND3X1 NAND3X1_482 ( .gnd(gnd), .vdd(vdd), .A(_2315_), .B(_343_), .C(_2321_), .Y(_2322_) );
NAND3X1 NAND3X1_483 ( .gnd(gnd), .vdd(vdd), .A(_2089_), .B(_2314_), .C(_2322_), .Y(_2323_) );
NAND3X1 NAND3X1_484 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_172_), .B(_343_), .C(_2321_), .Y(_2324_) );
OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_2313_), .B(_2311_), .C(_2315_), .Y(_2325_) );
NAND3X1 NAND3X1_485 ( .gnd(gnd), .vdd(vdd), .A(_1662_), .B(_2325_), .C(_2324_), .Y(_2326_) );
AOI21X1 AOI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_2323_), .B(_2326_), .C(_2088_), .Y(_2327_) );
INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .Y(_2328_) );
AOI21X1 AOI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_2328_), .B(_1545_), .C(_1664_), .Y(_2330_) );
AOI21X1 AOI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_2325_), .B(_2324_), .C(_1662_), .Y(_2331_) );
AOI21X1 AOI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_2314_), .B(_2322_), .C(_2089_), .Y(_2332_) );
NOR3X1 NOR3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_2331_), .B(_2332_), .C(_2330_), .Y(_2333_) );
OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_2333_), .B(_2327_), .C(_2482_), .Y(_2334_) );
OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_2332_), .B(_2331_), .C(_2330_), .Y(_2335_) );
NAND3X1 NAND3X1_486 ( .gnd(gnd), .vdd(vdd), .A(_2088_), .B(_2323_), .C(_2326_), .Y(_2336_) );
NAND3X1 NAND3X1_487 ( .gnd(gnd), .vdd(vdd), .A(_2285_), .B(_2336_), .C(_2335_), .Y(_2337_) );
NAND3X1 NAND3X1_488 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_2337_), .C(_2334_), .Y(_2338_) );
NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_188_), .B(_2338_), .Y(_2339_) );
INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_188_), .Y(_2341_) );
NAND3X1 NAND3X1_489 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_2336_), .C(_2335_), .Y(_2342_) );
OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_2333_), .B(_2327_), .C(_2285_), .Y(_2343_) );
NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_2342_), .B(_2343_), .Y(_2344_) );
NAND3X1 NAND3X1_490 ( .gnd(gnd), .vdd(vdd), .A(_2341_), .B(_362_), .C(_2344_), .Y(_2345_) );
NAND3X1 NAND3X1_491 ( .gnd(gnd), .vdd(vdd), .A(_2085_), .B(_2339_), .C(_2345_), .Y(_2346_) );
NAND3X1 NAND3X1_492 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_188_), .B(_362_), .C(_2344_), .Y(_2347_) );
NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_2341_), .B(_2338_), .Y(_2348_) );
NAND3X1 NAND3X1_493 ( .gnd(gnd), .vdd(vdd), .A(_1672_), .B(_2347_), .C(_2348_), .Y(_2349_) );
AOI21X1 AOI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_2346_), .B(_2349_), .C(_2084_), .Y(_2350_) );
INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(_1675_), .Y(_2352_) );
AOI21X1 AOI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1542_), .B(_2352_), .C(_1674_), .Y(_2353_) );
AOI21X1 AOI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_2347_), .B(_2348_), .C(_1672_), .Y(_2354_) );
AOI21X1 AOI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .B(_2345_), .C(_2085_), .Y(_2355_) );
NOR3X1 NOR3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_2354_), .B(_2355_), .C(_2353_), .Y(_2356_) );
OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_2356_), .B(_2350_), .C(_2318_), .Y(_2357_) );
OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_2355_), .B(_2354_), .C(_2353_), .Y(_2358_) );
NAND3X1 NAND3X1_494 ( .gnd(gnd), .vdd(vdd), .A(_2084_), .B(_2346_), .C(_2349_), .Y(_2359_) );
NAND3X1 NAND3X1_495 ( .gnd(gnd), .vdd(vdd), .A(_2449_), .B(_2359_), .C(_2358_), .Y(_2360_) );
NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_2360_), .B(_2357_), .Y(_2361_) );
NAND3X1 NAND3X1_496 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_204_), .B(_389_), .C(_2361_), .Y(_2363_) );
INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_204_), .Y(_2364_) );
AOI21X1 AOI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_2359_), .B(_2358_), .C(_2318_), .Y(_2365_) );
NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_2359_), .B(_2358_), .Y(_2366_) );
OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_2366_), .B(_2449_), .C(_389_), .Y(_2367_) );
OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_2367_), .B(_2365_), .C(_2364_), .Y(_2368_) );
AOI21X1 AOI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_2368_), .B(_2363_), .C(_1683_), .Y(_2369_) );
OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2367_), .B(_2365_), .C(module_0_W_204_), .Y(_2370_) );
NAND3X1 NAND3X1_497 ( .gnd(gnd), .vdd(vdd), .A(_2364_), .B(_389_), .C(_2361_), .Y(_2371_) );
AOI21X1 AOI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2370_), .B(_2371_), .C(_1682_), .Y(_2372_) );
OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_2372_), .B(_2369_), .C(_2083_), .Y(_2374_) );
AOI21X1 AOI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .B(_1683_), .C(_1445_), .Y(_2375_) );
OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_2375_), .B(_1540_), .C(_1684_), .Y(_2376_) );
NAND3X1 NAND3X1_498 ( .gnd(gnd), .vdd(vdd), .A(_1682_), .B(_2370_), .C(_2371_), .Y(_2377_) );
NAND3X1 NAND3X1_499 ( .gnd(gnd), .vdd(vdd), .A(_1683_), .B(_2368_), .C(_2363_), .Y(_2378_) );
NAND3X1 NAND3X1_500 ( .gnd(gnd), .vdd(vdd), .A(_2377_), .B(_2378_), .C(_2376_), .Y(_2379_) );
NAND3X1 NAND3X1_501 ( .gnd(gnd), .vdd(vdd), .A(_2428_), .B(_2379_), .C(_2374_), .Y(_2380_) );
AOI21X1 AOI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_2377_), .B(_2378_), .C(_2376_), .Y(_2381_) );
NOR3X1 NOR3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_2369_), .B(_2083_), .C(_2372_), .Y(_2382_) );
OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_2382_), .B(_2381_), .C(_2351_), .Y(_2383_) );
NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_2380_), .B(_2383_), .Y(_2385_) );
NAND3X1 NAND3X1_502 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_220_), .B(_410_), .C(_2385_), .Y(_2386_) );
INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_220_), .Y(_2387_) );
AOI21X1 AOI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_2379_), .B(_2374_), .C(_2351_), .Y(_2388_) );
NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_2379_), .B(_2374_), .Y(_2389_) );
OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .B(_2428_), .C(_410_), .Y(_2390_) );
OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2390_), .B(_2388_), .C(_2387_), .Y(_2391_) );
AOI21X1 AOI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_2391_), .B(_2386_), .C(_1696_), .Y(_2392_) );
OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_2390_), .B(_2388_), .C(module_0_W_220_), .Y(_2393_) );
NAND3X1 NAND3X1_503 ( .gnd(gnd), .vdd(vdd), .A(_2387_), .B(_410_), .C(_2385_), .Y(_2394_) );
AOI21X1 AOI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_2393_), .B(_2394_), .C(_1693_), .Y(_2396_) );
OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_2392_), .B(_2396_), .C(_2081_), .Y(_2397_) );
AOI21X1 AOI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_1479_), .B(_1487_), .C(_1489_), .Y(_2398_) );
NAND3X1 NAND3X1_504 ( .gnd(gnd), .vdd(vdd), .A(_1482_), .B(_1696_), .C(_1695_), .Y(_2399_) );
OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .B(_1697_), .C(_2399_), .Y(_2400_) );
NAND3X1 NAND3X1_505 ( .gnd(gnd), .vdd(vdd), .A(_1693_), .B(_2393_), .C(_2394_), .Y(_2401_) );
NAND3X1 NAND3X1_506 ( .gnd(gnd), .vdd(vdd), .A(_1696_), .B(_2391_), .C(_2386_), .Y(_2402_) );
NAND3X1 NAND3X1_507 ( .gnd(gnd), .vdd(vdd), .A(_2400_), .B(_2401_), .C(_2402_), .Y(_2403_) );
AOI21X1 AOI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_2403_), .B(_2397_), .C(_2384_), .Y(_2404_) );
NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_2403_), .B(_2397_), .Y(_2405_) );
OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_2405_), .B(_2395_), .C(_436_), .Y(_2407_) );
OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_2407_), .B(_2404_), .C(module_0_W_236_), .Y(_2408_) );
INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_236_), .Y(_2409_) );
NAND3X1 NAND3X1_508 ( .gnd(gnd), .vdd(vdd), .A(_2395_), .B(_2403_), .C(_2397_), .Y(_2410_) );
AOI21X1 AOI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_2401_), .B(_2402_), .C(_2400_), .Y(_2411_) );
NOR3X1 NOR3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_2392_), .B(_2081_), .C(_2396_), .Y(_2412_) );
OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_2412_), .B(_2411_), .C(_2384_), .Y(_2413_) );
NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_2410_), .B(_2413_), .Y(_2414_) );
NAND3X1 NAND3X1_509 ( .gnd(gnd), .vdd(vdd), .A(_2409_), .B(_436_), .C(_2414_), .Y(_2415_) );
NAND3X1 NAND3X1_510 ( .gnd(gnd), .vdd(vdd), .A(_2079_), .B(_2408_), .C(_2415_), .Y(_2416_) );
NAND3X1 NAND3X1_511 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_236_), .B(_436_), .C(_2414_), .Y(_2418_) );
OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_2407_), .B(_2404_), .C(_2409_), .Y(_2419_) );
NAND3X1 NAND3X1_512 ( .gnd(gnd), .vdd(vdd), .A(_1703_), .B(_2419_), .C(_2418_), .Y(_2420_) );
AOI21X1 AOI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_2416_), .B(_2420_), .C(_2078_), .Y(_2421_) );
INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(_1706_), .Y(_2422_) );
AOI21X1 AOI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_1709_), .B(_2422_), .C(_1705_), .Y(_2423_) );
NAND3X1 NAND3X1_513 ( .gnd(gnd), .vdd(vdd), .A(_2079_), .B(_2419_), .C(_2418_), .Y(_2424_) );
NAND3X1 NAND3X1_514 ( .gnd(gnd), .vdd(vdd), .A(_1703_), .B(_2408_), .C(_2415_), .Y(_2425_) );
AOI21X1 AOI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_2424_), .B(_2425_), .C(_2423_), .Y(_2426_) );
OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_2426_), .B(_2421_), .C(_3629_), .Y(_2427_) );
AOI21X1 AOI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_2419_), .B(_2418_), .C(_1703_), .Y(_2429_) );
AOI21X1 AOI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2408_), .B(_2415_), .C(_2079_), .Y(_2430_) );
OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_2429_), .B(_2430_), .C(_2423_), .Y(_2431_) );
NAND3X1 NAND3X1_515 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .B(_2416_), .C(_2420_), .Y(_2432_) );
NAND3X1 NAND3X1_516 ( .gnd(gnd), .vdd(vdd), .A(_3630_), .B(_2432_), .C(_2431_), .Y(_2433_) );
NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_2433_), .B(_2427_), .Y(_2434_) );
NAND3X1 NAND3X1_517 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_252_), .B(_460_), .C(_2434_), .Y(_2435_) );
INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_252_), .Y(_2436_) );
AOI21X1 AOI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_2432_), .B(_2431_), .C(_3629_), .Y(_2437_) );
NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2432_), .B(_2431_), .Y(_2438_) );
OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_2438_), .B(_3630_), .C(_460_), .Y(_2440_) );
OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_2440_), .B(_2437_), .C(_2436_), .Y(_2441_) );
AOI21X1 AOI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_2441_), .B(_2435_), .C(_2070_), .Y(_2442_) );
INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(_2442_), .Y(_2443_) );
NAND3X1 NAND3X1_518 ( .gnd(gnd), .vdd(vdd), .A(_2070_), .B(_2441_), .C(_2435_), .Y(_2444_) );
NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_2444_), .B(_2443_), .Y(_2445_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_2445_), .B(_2077_), .Y(module_0_H_20_) );
OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_2442_), .B(_2077_), .C(_2444_), .Y(_2446_) );
NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_2434_), .Y(_2447_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_252_), .B(_2447_), .Y(_2448_) );
AOI21X1 AOI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .B(_2420_), .C(_2429_), .Y(_2450_) );
INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_237_), .Y(_2451_) );
OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_2396_), .B(_2081_), .C(_2401_), .Y(_2452_) );
INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(_2393_), .Y(_2453_) );
AOI21X1 AOI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_2378_), .B(_2376_), .C(_2369_), .Y(_2454_) );
INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_205_), .Y(_2455_) );
OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_2353_), .B(_2355_), .C(_2346_), .Y(_2456_) );
INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .Y(_2457_) );
AOI21X1 AOI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_2088_), .B(_2326_), .C(_2331_), .Y(_2458_) );
INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_173_), .Y(_2459_) );
INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(_3400_), .Y(_2461_) );
AOI21X1 AOI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_2306_), .B(_2309_), .C(_2300_), .Y(_2462_) );
INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_157_), .Y(_2463_) );
INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(_3316_), .Y(_2464_) );
AOI21X1 AOI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_2092_), .B(_2287_), .C(_2279_), .Y(_2465_) );
INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_141_), .Y(_2466_) );
OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_2260_), .B(_2095_), .C(_2264_), .Y(_2467_) );
INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf3_), .Y(_2468_) );
AOI21X1 AOI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_2239_), .B(_2100_), .C(_2244_), .Y(_2469_) );
INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(_2237_), .Y(_2470_) );
INVX1 INVX1_264 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf4_), .Y(_2472_) );
AOI21X1 AOI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_2216_), .B(_2104_), .C(_2221_), .Y(_2473_) );
INVX1 INVX1_265 ( .gnd(gnd), .vdd(vdd), .A(_2214_), .Y(_2474_) );
INVX1 INVX1_266 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf4_), .Y(_2475_) );
AOI21X1 AOI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2199_), .B(_2196_), .C(_2190_), .Y(_2476_) );
INVX1 INVX1_267 ( .gnd(gnd), .vdd(vdd), .A(_2185_), .Y(_2477_) );
INVX1 INVX1_268 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf4_), .Y(_2478_) );
OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .B(_2172_), .C(_2176_), .Y(_2479_) );
INVX1 INVX1_269 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf4_), .Y(_2480_) );
AOI21X1 AOI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2151_), .B(_2116_), .C(_2156_), .Y(_2481_) );
INVX1 INVX1_270 ( .gnd(gnd), .vdd(vdd), .A(_2149_), .Y(_2483_) );
INVX1 INVX1_271 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf3_), .Y(_2484_) );
OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_2135_), .B(_2134_), .C(_2130_), .Y(_2485_) );
INVX1 INVX1_272 ( .gnd(gnd), .vdd(vdd), .A(_2125_), .Y(_2486_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_12_), .B(module_0_W_13_), .Y(_2487_) );
INVX1 INVX1_273 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .Y(_2488_) );
OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .B(_2779_), .C(module_0_W_9_), .Y(_2489_) );
NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_629_), .Y(_2490_) );
NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_2489_), .B(_2490_), .Y(_2491_) );
NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_2488_), .B(_2491_), .Y(_2492_) );
NAND3X1 NAND3X1_519 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .B(_2489_), .C(_2490_), .Y(_2494_) );
AOI21X1 AOI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2494_), .B(_2492_), .C(module_0_W_29_), .Y(_2495_) );
INVX1 INVX1_274 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_29_), .Y(_2496_) );
NAND2X1 NAND2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .B(_2491_), .Y(_2497_) );
NAND3X1 NAND3X1_520 ( .gnd(gnd), .vdd(vdd), .A(_2488_), .B(_2489_), .C(_2490_), .Y(_2498_) );
AOI21X1 AOI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_2498_), .B(_2497_), .C(_2496_), .Y(_2499_) );
OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_2499_), .B(_2495_), .C(_2486_), .Y(_2500_) );
NAND3X1 NAND3X1_521 ( .gnd(gnd), .vdd(vdd), .A(_2496_), .B(_2498_), .C(_2497_), .Y(_2501_) );
NAND3X1 NAND3X1_522 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_29_), .B(_2494_), .C(_2492_), .Y(_2502_) );
NAND3X1 NAND3X1_523 ( .gnd(gnd), .vdd(vdd), .A(_2125_), .B(_2502_), .C(_2501_), .Y(_2503_) );
NAND3X1 NAND3X1_524 ( .gnd(gnd), .vdd(vdd), .A(_2500_), .B(_2503_), .C(_2485_), .Y(_2505_) );
AOI21X1 AOI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_2128_), .B(_2121_), .C(_2129_), .Y(_2506_) );
AOI21X1 AOI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_2502_), .B(_2501_), .C(_2125_), .Y(_2507_) );
NOR3X1 NOR3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_2495_), .B(_2486_), .C(_2499_), .Y(_2508_) );
OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_2508_), .B(_2507_), .C(_2506_), .Y(_2509_) );
XNOR2X1 XNOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_492_), .B(_2855_), .Y(_2510_) );
INVX1 INVX1_275 ( .gnd(gnd), .vdd(vdd), .A(_2510_), .Y(_2511_) );
NAND3X1 NAND3X1_525 ( .gnd(gnd), .vdd(vdd), .A(_2509_), .B(_2511_), .C(_2505_), .Y(_2512_) );
NOR3X1 NOR3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_2506_), .B(_2507_), .C(_2508_), .Y(_2513_) );
AOI21X1 AOI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_2500_), .B(_2503_), .C(_2485_), .Y(_2514_) );
OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .B(_2514_), .C(_2510_), .Y(_2516_) );
NAND3X1 NAND3X1_526 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .B(_2512_), .C(_2516_), .Y(_2517_) );
NAND3X1 NAND3X1_527 ( .gnd(gnd), .vdd(vdd), .A(_2509_), .B(_2510_), .C(_2505_), .Y(_2518_) );
OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .B(_2514_), .C(_2511_), .Y(_2519_) );
NAND3X1 NAND3X1_528 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf2_), .B(_2518_), .C(_2519_), .Y(_2520_) );
NAND3X1 NAND3X1_529 ( .gnd(gnd), .vdd(vdd), .A(_2483_), .B(_2517_), .C(_2520_), .Y(_2521_) );
AOI21X1 AOI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_2518_), .B(_2519_), .C(bloque_datos_13_bF_buf1_), .Y(_2522_) );
AOI21X1 AOI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_2512_), .B(_2516_), .C(_2484_), .Y(_2523_) );
OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_2522_), .B(_2523_), .C(_2149_), .Y(_2524_) );
NAND3X1 NAND3X1_530 ( .gnd(gnd), .vdd(vdd), .A(_2521_), .B(_2524_), .C(_2481_), .Y(_2525_) );
OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_2157_), .B(_2155_), .C(_2147_), .Y(_2527_) );
NAND3X1 NAND3X1_531 ( .gnd(gnd), .vdd(vdd), .A(_2149_), .B(_2517_), .C(_2520_), .Y(_2528_) );
OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_2522_), .B(_2523_), .C(_2483_), .Y(_2529_) );
NAND3X1 NAND3X1_532 ( .gnd(gnd), .vdd(vdd), .A(_2528_), .B(_2529_), .C(_2527_), .Y(_2530_) );
XNOR2X1 XNOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(_2899_), .Y(_2531_) );
INVX1 INVX1_276 ( .gnd(gnd), .vdd(vdd), .A(_2531_), .Y(_2532_) );
NAND3X1 NAND3X1_533 ( .gnd(gnd), .vdd(vdd), .A(_2530_), .B(_2532_), .C(_2525_), .Y(_2533_) );
AOI21X1 AOI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_2528_), .B(_2529_), .C(_2527_), .Y(_2534_) );
AOI21X1 AOI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_2521_), .B(_2524_), .C(_2481_), .Y(_2535_) );
OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_2535_), .B(_2534_), .C(_2531_), .Y(_2536_) );
NAND3X1 NAND3X1_534 ( .gnd(gnd), .vdd(vdd), .A(_2480_), .B(_2533_), .C(_2536_), .Y(_2538_) );
NOR3X1 NOR3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_2534_), .B(_2531_), .C(_2535_), .Y(_2539_) );
AOI21X1 AOI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_2530_), .B(_2525_), .C(_2532_), .Y(_2540_) );
OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_2539_), .B(_2540_), .C(bloque_datos_29_bF_buf3_), .Y(_2541_) );
NAND3X1 NAND3X1_535 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(_2538_), .C(_2541_), .Y(_2542_) );
INVX1 INVX1_277 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .Y(_2543_) );
NOR3X1 NOR3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_2540_), .B(bloque_datos_29_bF_buf2_), .C(_2539_), .Y(_2544_) );
AOI21X1 AOI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_2533_), .B(_2536_), .C(_2480_), .Y(_2545_) );
OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_2544_), .B(_2545_), .C(_2543_), .Y(_2546_) );
AOI21X1 AOI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_2542_), .B(_2546_), .C(_2479_), .Y(_2547_) );
AOI21X1 AOI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_2177_), .B(_2174_), .C(_2168_), .Y(_2549_) );
NAND3X1 NAND3X1_536 ( .gnd(gnd), .vdd(vdd), .A(_2543_), .B(_2538_), .C(_2541_), .Y(_2550_) );
OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_2544_), .B(_2545_), .C(_2163_), .Y(_2551_) );
AOI21X1 AOI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2550_), .B(_2551_), .C(_2549_), .Y(_2552_) );
XNOR2X1 XNOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_2954_), .Y(_2553_) );
NOR3X1 NOR3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .B(_2553_), .C(_2547_), .Y(_2554_) );
NAND3X1 NAND3X1_537 ( .gnd(gnd), .vdd(vdd), .A(_2550_), .B(_2549_), .C(_2551_), .Y(_2555_) );
NAND3X1 NAND3X1_538 ( .gnd(gnd), .vdd(vdd), .A(_2479_), .B(_2542_), .C(_2546_), .Y(_2556_) );
INVX1 INVX1_278 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .Y(_2557_) );
AOI21X1 AOI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_2555_), .B(_2556_), .C(_2557_), .Y(_2558_) );
OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_2554_), .B(_2558_), .C(_2478_), .Y(_2560_) );
NAND3X1 NAND3X1_539 ( .gnd(gnd), .vdd(vdd), .A(_2557_), .B(_2555_), .C(_2556_), .Y(_2561_) );
OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .B(_2552_), .C(_2553_), .Y(_2562_) );
NAND3X1 NAND3X1_540 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf3_), .B(_2561_), .C(_2562_), .Y(_2563_) );
NAND3X1 NAND3X1_541 ( .gnd(gnd), .vdd(vdd), .A(_2477_), .B(_2563_), .C(_2560_), .Y(_2564_) );
AOI21X1 AOI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_2561_), .B(_2562_), .C(bloque_datos_45_bF_buf2_), .Y(_2565_) );
NOR3X1 NOR3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_2558_), .B(_2478_), .C(_2554_), .Y(_2566_) );
OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_2566_), .B(_2565_), .C(_2185_), .Y(_2567_) );
NAND3X1 NAND3X1_542 ( .gnd(gnd), .vdd(vdd), .A(_2564_), .B(_2567_), .C(_2476_), .Y(_2568_) );
OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_2107_), .B(_2193_), .C(_2198_), .Y(_2569_) );
NAND3X1 NAND3X1_543 ( .gnd(gnd), .vdd(vdd), .A(_2185_), .B(_2563_), .C(_2560_), .Y(_2571_) );
OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_2566_), .B(_2565_), .C(_2477_), .Y(_2572_) );
NAND3X1 NAND3X1_544 ( .gnd(gnd), .vdd(vdd), .A(_2571_), .B(_2569_), .C(_2572_), .Y(_2573_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_517_), .B(_3031_), .Y(_2574_) );
INVX1 INVX1_279 ( .gnd(gnd), .vdd(vdd), .A(_2574_), .Y(_2575_) );
NAND3X1 NAND3X1_545 ( .gnd(gnd), .vdd(vdd), .A(_2575_), .B(_2573_), .C(_2568_), .Y(_2576_) );
AOI21X1 AOI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_2571_), .B(_2572_), .C(_2569_), .Y(_2577_) );
AOI21X1 AOI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_2564_), .B(_2567_), .C(_2476_), .Y(_2578_) );
OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_2578_), .B(_2577_), .C(_2574_), .Y(_2579_) );
NAND3X1 NAND3X1_546 ( .gnd(gnd), .vdd(vdd), .A(_2475_), .B(_2576_), .C(_2579_), .Y(_2580_) );
NAND3X1 NAND3X1_547 ( .gnd(gnd), .vdd(vdd), .A(_2574_), .B(_2573_), .C(_2568_), .Y(_2582_) );
OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_2578_), .B(_2577_), .C(_2575_), .Y(_2583_) );
NAND3X1 NAND3X1_548 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf3_), .B(_2582_), .C(_2583_), .Y(_2584_) );
NAND3X1 NAND3X1_549 ( .gnd(gnd), .vdd(vdd), .A(_2474_), .B(_2580_), .C(_2584_), .Y(_2585_) );
AOI21X1 AOI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2582_), .B(_2583_), .C(bloque_datos_61_bF_buf2_), .Y(_2586_) );
AOI21X1 AOI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_2576_), .B(_2579_), .C(_2475_), .Y(_2587_) );
OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2586_), .B(_2587_), .C(_2214_), .Y(_2588_) );
NAND3X1 NAND3X1_550 ( .gnd(gnd), .vdd(vdd), .A(_2585_), .B(_2588_), .C(_2473_), .Y(_2589_) );
OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2220_), .B(_2222_), .C(_2212_), .Y(_2590_) );
NAND3X1 NAND3X1_551 ( .gnd(gnd), .vdd(vdd), .A(_2214_), .B(_2580_), .C(_2584_), .Y(_2591_) );
OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_2586_), .B(_2587_), .C(_2474_), .Y(_2593_) );
NAND3X1 NAND3X1_552 ( .gnd(gnd), .vdd(vdd), .A(_2591_), .B(_2590_), .C(_2593_), .Y(_2594_) );
XNOR2X1 XNOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_3097_), .Y(_2595_) );
INVX1 INVX1_280 ( .gnd(gnd), .vdd(vdd), .A(_2595_), .Y(_2596_) );
NAND3X1 NAND3X1_553 ( .gnd(gnd), .vdd(vdd), .A(_2596_), .B(_2594_), .C(_2589_), .Y(_2597_) );
AOI21X1 AOI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_2591_), .B(_2593_), .C(_2590_), .Y(_2598_) );
AOI21X1 AOI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_2585_), .B(_2588_), .C(_2473_), .Y(_2599_) );
OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_2598_), .B(_2599_), .C(_2595_), .Y(_2600_) );
NAND3X1 NAND3X1_554 ( .gnd(gnd), .vdd(vdd), .A(_2472_), .B(_2597_), .C(_2600_), .Y(_2601_) );
NAND3X1 NAND3X1_555 ( .gnd(gnd), .vdd(vdd), .A(_2595_), .B(_2594_), .C(_2589_), .Y(_2602_) );
OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_2598_), .B(_2599_), .C(_2596_), .Y(_2604_) );
NAND3X1 NAND3X1_556 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf3_), .B(_2602_), .C(_2604_), .Y(_2605_) );
NAND3X1 NAND3X1_557 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .B(_2601_), .C(_2605_), .Y(_2606_) );
AOI21X1 AOI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_2602_), .B(_2604_), .C(bloque_datos_77_bF_buf2_), .Y(_2607_) );
AOI21X1 AOI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_2597_), .B(_2600_), .C(_2472_), .Y(_2608_) );
OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_2607_), .B(_2608_), .C(_2237_), .Y(_2609_) );
NAND3X1 NAND3X1_558 ( .gnd(gnd), .vdd(vdd), .A(_2606_), .B(_2609_), .C(_2469_), .Y(_2610_) );
OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2245_), .B(_2243_), .C(_2235_), .Y(_2611_) );
NAND3X1 NAND3X1_559 ( .gnd(gnd), .vdd(vdd), .A(_2237_), .B(_2601_), .C(_2605_), .Y(_2612_) );
OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_2607_), .B(_2608_), .C(_2470_), .Y(_2613_) );
NAND3X1 NAND3X1_560 ( .gnd(gnd), .vdd(vdd), .A(_2612_), .B(_2611_), .C(_2613_), .Y(_2615_) );
XNOR2X1 XNOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_3141_), .Y(_2616_) );
INVX1 INVX1_281 ( .gnd(gnd), .vdd(vdd), .A(_2616_), .Y(_2617_) );
NAND3X1 NAND3X1_561 ( .gnd(gnd), .vdd(vdd), .A(_2617_), .B(_2615_), .C(_2610_), .Y(_2618_) );
AOI21X1 AOI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_2612_), .B(_2613_), .C(_2611_), .Y(_2619_) );
AOI21X1 AOI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_2606_), .B(_2609_), .C(_2469_), .Y(_2620_) );
OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_2619_), .B(_2620_), .C(_2616_), .Y(_2621_) );
NAND3X1 NAND3X1_562 ( .gnd(gnd), .vdd(vdd), .A(_2468_), .B(_2618_), .C(_2621_), .Y(_2622_) );
NOR3X1 NOR3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_2619_), .B(_2616_), .C(_2620_), .Y(_2623_) );
AOI21X1 AOI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_2615_), .B(_2610_), .C(_2617_), .Y(_2624_) );
OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_2623_), .B(_2624_), .C(bloque_datos_93_bF_buf2_), .Y(_2626_) );
NAND3X1 NAND3X1_563 ( .gnd(gnd), .vdd(vdd), .A(_2253_), .B(_2622_), .C(_2626_), .Y(_2627_) );
INVX1 INVX1_282 ( .gnd(gnd), .vdd(vdd), .A(_2253_), .Y(_2628_) );
NOR3X1 NOR3X1_61 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf1_), .B(_2624_), .C(_2623_), .Y(_2629_) );
AOI21X1 AOI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_2618_), .B(_2621_), .C(_2468_), .Y(_2630_) );
OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_2629_), .B(_2630_), .C(_2628_), .Y(_2631_) );
AOI21X1 AOI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_2627_), .B(_2631_), .C(_2467_), .Y(_2632_) );
AOI21X1 AOI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_2262_), .B(_2265_), .C(_2257_), .Y(_2633_) );
NAND3X1 NAND3X1_564 ( .gnd(gnd), .vdd(vdd), .A(_2628_), .B(_2622_), .C(_2626_), .Y(_2634_) );
OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_2629_), .B(_2630_), .C(_2253_), .Y(_2635_) );
AOI21X1 AOI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_2634_), .B(_2635_), .C(_2633_), .Y(_2637_) );
OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_2632_), .B(_2637_), .C(_3239_), .Y(_2638_) );
NAND3X1 NAND3X1_565 ( .gnd(gnd), .vdd(vdd), .A(_2633_), .B(_2634_), .C(_2635_), .Y(_2639_) );
NAND3X1 NAND3X1_566 ( .gnd(gnd), .vdd(vdd), .A(_2467_), .B(_2627_), .C(_2631_), .Y(_2640_) );
NAND3X1 NAND3X1_567 ( .gnd(gnd), .vdd(vdd), .A(_3250_), .B(_2639_), .C(_2640_), .Y(_2641_) );
NAND2X1 NAND2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_2641_), .B(_2638_), .Y(_2642_) );
NAND3X1 NAND3X1_568 ( .gnd(gnd), .vdd(vdd), .A(_2466_), .B(_535_), .C(_2642_), .Y(_2643_) );
OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_2632_), .B(_2637_), .C(_3250_), .Y(_2644_) );
NAND3X1 NAND3X1_569 ( .gnd(gnd), .vdd(vdd), .A(_3239_), .B(_2639_), .C(_2640_), .Y(_2645_) );
NAND3X1 NAND3X1_570 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_2645_), .C(_2644_), .Y(_2646_) );
NAND2X1 NAND2X1_326 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_141_), .B(_2646_), .Y(_2648_) );
AOI21X1 AOI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_2643_), .B(_2648_), .C(_2281_), .Y(_2649_) );
INVX1 INVX1_283 ( .gnd(gnd), .vdd(vdd), .A(_2281_), .Y(_2650_) );
NAND3X1 NAND3X1_571 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_141_), .B(_535_), .C(_2642_), .Y(_2651_) );
NAND2X1 NAND2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_2466_), .B(_2646_), .Y(_2652_) );
AOI21X1 AOI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_2651_), .B(_2652_), .C(_2650_), .Y(_2653_) );
OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_2649_), .B(_2653_), .C(_2465_), .Y(_2654_) );
OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_2093_), .B(_2283_), .C(_2286_), .Y(_2655_) );
NAND3X1 NAND3X1_572 ( .gnd(gnd), .vdd(vdd), .A(_2650_), .B(_2651_), .C(_2652_), .Y(_2656_) );
NAND3X1 NAND3X1_573 ( .gnd(gnd), .vdd(vdd), .A(_2281_), .B(_2643_), .C(_2648_), .Y(_2657_) );
NAND3X1 NAND3X1_574 ( .gnd(gnd), .vdd(vdd), .A(_2656_), .B(_2657_), .C(_2655_), .Y(_2659_) );
NAND3X1 NAND3X1_575 ( .gnd(gnd), .vdd(vdd), .A(_2464_), .B(_2659_), .C(_2654_), .Y(_2660_) );
AOI21X1 AOI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_2656_), .B(_2657_), .C(_2655_), .Y(_2661_) );
NOR3X1 NOR3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_2649_), .B(_2465_), .C(_2653_), .Y(_2662_) );
OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_2662_), .B(_2661_), .C(_3316_), .Y(_2663_) );
NAND2X1 NAND2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_2660_), .B(_2663_), .Y(_2664_) );
NAND3X1 NAND3X1_576 ( .gnd(gnd), .vdd(vdd), .A(_2463_), .B(_543_), .C(_2664_), .Y(_2665_) );
OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_2662_), .B(_2661_), .C(_2464_), .Y(_2666_) );
NAND3X1 NAND3X1_577 ( .gnd(gnd), .vdd(vdd), .A(_3316_), .B(_2659_), .C(_2654_), .Y(_2667_) );
NAND3X1 NAND3X1_578 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_2667_), .C(_2666_), .Y(_2668_) );
NAND2X1 NAND2X1_329 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_157_), .B(_2668_), .Y(_2670_) );
AOI21X1 AOI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_2665_), .B(_2670_), .C(_2301_), .Y(_2671_) );
INVX1 INVX1_284 ( .gnd(gnd), .vdd(vdd), .A(_2301_), .Y(_2672_) );
NAND3X1 NAND3X1_579 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_157_), .B(_543_), .C(_2664_), .Y(_2673_) );
NAND2X1 NAND2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_2463_), .B(_2668_), .Y(_2674_) );
AOI21X1 AOI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_2673_), .B(_2674_), .C(_2672_), .Y(_2675_) );
OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_2671_), .B(_2675_), .C(_2462_), .Y(_2676_) );
OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_2303_), .B(_2091_), .C(_2308_), .Y(_2677_) );
NAND3X1 NAND3X1_580 ( .gnd(gnd), .vdd(vdd), .A(_2672_), .B(_2673_), .C(_2674_), .Y(_2678_) );
NAND3X1 NAND3X1_581 ( .gnd(gnd), .vdd(vdd), .A(_2301_), .B(_2665_), .C(_2670_), .Y(_2679_) );
NAND3X1 NAND3X1_582 ( .gnd(gnd), .vdd(vdd), .A(_2678_), .B(_2679_), .C(_2677_), .Y(_2681_) );
NAND3X1 NAND3X1_583 ( .gnd(gnd), .vdd(vdd), .A(_2461_), .B(_2681_), .C(_2676_), .Y(_2682_) );
AOI21X1 AOI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_2678_), .B(_2679_), .C(_2677_), .Y(_2683_) );
NOR3X1 NOR3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_2671_), .B(_2462_), .C(_2675_), .Y(_2684_) );
OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_2684_), .B(_2683_), .C(_3400_), .Y(_2685_) );
NAND2X1 NAND2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2682_), .B(_2685_), .Y(_2686_) );
NAND3X1 NAND3X1_584 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .B(_551_), .C(_2686_), .Y(_2687_) );
OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_2684_), .B(_2683_), .C(_2461_), .Y(_2688_) );
NAND3X1 NAND3X1_585 ( .gnd(gnd), .vdd(vdd), .A(_3400_), .B(_2681_), .C(_2676_), .Y(_2689_) );
NAND3X1 NAND3X1_586 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_2689_), .C(_2688_), .Y(_2690_) );
NAND2X1 NAND2X1_332 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_173_), .B(_2690_), .Y(_2692_) );
AOI21X1 AOI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_2687_), .B(_2692_), .C(_2314_), .Y(_2693_) );
INVX1 INVX1_285 ( .gnd(gnd), .vdd(vdd), .A(_2314_), .Y(_2694_) );
NAND3X1 NAND3X1_587 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_173_), .B(_551_), .C(_2686_), .Y(_2695_) );
NAND2X1 NAND2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .B(_2690_), .Y(_2696_) );
AOI21X1 AOI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_2695_), .B(_2696_), .C(_2694_), .Y(_2697_) );
OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_2693_), .B(_2697_), .C(_2458_), .Y(_2698_) );
OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_2330_), .B(_2332_), .C(_2323_), .Y(_2699_) );
NAND3X1 NAND3X1_588 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .B(_2695_), .C(_2696_), .Y(_2700_) );
NAND3X1 NAND3X1_589 ( .gnd(gnd), .vdd(vdd), .A(_2314_), .B(_2687_), .C(_2692_), .Y(_2701_) );
NAND3X1 NAND3X1_590 ( .gnd(gnd), .vdd(vdd), .A(_2700_), .B(_2701_), .C(_2699_), .Y(_2703_) );
NAND3X1 NAND3X1_591 ( .gnd(gnd), .vdd(vdd), .A(_3409_), .B(_2703_), .C(_2698_), .Y(_2704_) );
AOI21X1 AOI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_2700_), .B(_2701_), .C(_2699_), .Y(_2705_) );
NOR3X1 NOR3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_2693_), .B(_2458_), .C(_2697_), .Y(_2706_) );
OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_2706_), .B(_2705_), .C(_3408_), .Y(_2707_) );
NAND2X1 NAND2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_2704_), .B(_2707_), .Y(_2708_) );
NAND3X1 NAND3X1_592 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_189_), .B(_559_), .C(_2708_), .Y(_2709_) );
INVX1 INVX1_286 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_189_), .Y(_2710_) );
OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_2706_), .B(_2705_), .C(_3409_), .Y(_2711_) );
NAND3X1 NAND3X1_593 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .B(_2703_), .C(_2698_), .Y(_2712_) );
NAND3X1 NAND3X1_594 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_2712_), .C(_2711_), .Y(_2714_) );
NAND2X1 NAND2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_2710_), .B(_2714_), .Y(_2715_) );
NAND3X1 NAND3X1_595 ( .gnd(gnd), .vdd(vdd), .A(_2457_), .B(_2709_), .C(_2715_), .Y(_2716_) );
NAND3X1 NAND3X1_596 ( .gnd(gnd), .vdd(vdd), .A(_2710_), .B(_559_), .C(_2708_), .Y(_2717_) );
NAND2X1 NAND2X1_336 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_189_), .B(_2714_), .Y(_2718_) );
NAND3X1 NAND3X1_597 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .B(_2717_), .C(_2718_), .Y(_2719_) );
AOI21X1 AOI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_2716_), .B(_2719_), .C(_2456_), .Y(_2720_) );
AOI21X1 AOI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_2084_), .B(_2349_), .C(_2354_), .Y(_2721_) );
AOI21X1 AOI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_2717_), .B(_2718_), .C(_2339_), .Y(_2722_) );
AOI21X1 AOI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_2709_), .B(_2715_), .C(_2457_), .Y(_2723_) );
NOR3X1 NOR3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_2722_), .B(_2721_), .C(_2723_), .Y(_2725_) );
OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_2725_), .B(_2720_), .C(_3417_), .Y(_2726_) );
INVX1 INVX1_287 ( .gnd(gnd), .vdd(vdd), .A(_3417_), .Y(_2727_) );
OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_2722_), .B(_2723_), .C(_2721_), .Y(_2728_) );
NAND3X1 NAND3X1_598 ( .gnd(gnd), .vdd(vdd), .A(_2716_), .B(_2719_), .C(_2456_), .Y(_2729_) );
NAND3X1 NAND3X1_599 ( .gnd(gnd), .vdd(vdd), .A(_2727_), .B(_2728_), .C(_2729_), .Y(_2730_) );
NAND2X1 NAND2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .B(_2726_), .Y(_2731_) );
NAND3X1 NAND3X1_600 ( .gnd(gnd), .vdd(vdd), .A(_2455_), .B(_567_), .C(_2731_), .Y(_2732_) );
OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_2725_), .B(_2720_), .C(_2727_), .Y(_2733_) );
NAND3X1 NAND3X1_601 ( .gnd(gnd), .vdd(vdd), .A(_3417_), .B(_2728_), .C(_2729_), .Y(_2734_) );
NAND3X1 NAND3X1_602 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_2734_), .C(_2733_), .Y(_2736_) );
NAND2X1 NAND2X1_338 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_205_), .B(_2736_), .Y(_2737_) );
AOI21X1 AOI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .B(_2737_), .C(_2370_), .Y(_2738_) );
INVX1 INVX1_288 ( .gnd(gnd), .vdd(vdd), .A(_2370_), .Y(_2739_) );
NAND3X1 NAND3X1_603 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_205_), .B(_567_), .C(_2731_), .Y(_2740_) );
NAND2X1 NAND2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_2455_), .B(_2736_), .Y(_2741_) );
AOI21X1 AOI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_2740_), .B(_2741_), .C(_2739_), .Y(_2742_) );
OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_2738_), .B(_2742_), .C(_2454_), .Y(_2743_) );
OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_2372_), .B(_2083_), .C(_2377_), .Y(_2744_) );
NAND3X1 NAND3X1_604 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2740_), .C(_2741_), .Y(_2745_) );
NAND3X1 NAND3X1_605 ( .gnd(gnd), .vdd(vdd), .A(_2370_), .B(_2732_), .C(_2737_), .Y(_2747_) );
NAND3X1 NAND3X1_606 ( .gnd(gnd), .vdd(vdd), .A(_2745_), .B(_2747_), .C(_2744_), .Y(_2748_) );
NAND3X1 NAND3X1_607 ( .gnd(gnd), .vdd(vdd), .A(_3425_), .B(_2748_), .C(_2743_), .Y(_2749_) );
NAND2X1 NAND2X1_340 ( .gnd(gnd), .vdd(vdd), .A(_2748_), .B(_2743_), .Y(_2750_) );
AOI21X1 AOI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_3426_), .B(_2750_), .C(_576_), .Y(_2751_) );
NAND3X1 NAND3X1_608 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_221_), .B(_2749_), .C(_2751_), .Y(_2752_) );
INVX1 INVX1_289 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_221_), .Y(_2753_) );
AOI21X1 AOI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_2745_), .B(_2747_), .C(_2744_), .Y(_2754_) );
NOR3X1 NOR3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_2454_), .B(_2738_), .C(_2742_), .Y(_2755_) );
OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_2755_), .B(_2754_), .C(_3426_), .Y(_2756_) );
NAND3X1 NAND3X1_609 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_2749_), .C(_2756_), .Y(_2758_) );
NAND2X1 NAND2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2753_), .B(_2758_), .Y(_2759_) );
NAND3X1 NAND3X1_610 ( .gnd(gnd), .vdd(vdd), .A(_2453_), .B(_2752_), .C(_2759_), .Y(_2760_) );
NAND3X1 NAND3X1_611 ( .gnd(gnd), .vdd(vdd), .A(_2753_), .B(_2749_), .C(_2751_), .Y(_2761_) );
NAND2X1 NAND2X1_342 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_221_), .B(_2758_), .Y(_2762_) );
NAND3X1 NAND3X1_612 ( .gnd(gnd), .vdd(vdd), .A(_2393_), .B(_2761_), .C(_2762_), .Y(_2763_) );
AOI21X1 AOI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_2760_), .B(_2763_), .C(_2452_), .Y(_2764_) );
AOI21X1 AOI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_2400_), .B(_2402_), .C(_2392_), .Y(_2765_) );
AOI21X1 AOI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_2761_), .B(_2762_), .C(_2393_), .Y(_2766_) );
AOI21X1 AOI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_2752_), .B(_2759_), .C(_2453_), .Y(_2767_) );
NOR3X1 NOR3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_2766_), .B(_2765_), .C(_2767_), .Y(_2769_) );
OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_2769_), .B(_2764_), .C(_3434_), .Y(_2770_) );
INVX1 INVX1_290 ( .gnd(gnd), .vdd(vdd), .A(_3434_), .Y(_2771_) );
OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_2766_), .B(_2767_), .C(_2765_), .Y(_2772_) );
NAND3X1 NAND3X1_613 ( .gnd(gnd), .vdd(vdd), .A(_2760_), .B(_2763_), .C(_2452_), .Y(_2773_) );
NAND3X1 NAND3X1_614 ( .gnd(gnd), .vdd(vdd), .A(_2771_), .B(_2773_), .C(_2772_), .Y(_2774_) );
NAND2X1 NAND2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2774_), .B(_2770_), .Y(_2775_) );
NAND3X1 NAND3X1_615 ( .gnd(gnd), .vdd(vdd), .A(_2451_), .B(_583_), .C(_2775_), .Y(_2776_) );
OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_2769_), .B(_2764_), .C(_2771_), .Y(_2777_) );
NAND3X1 NAND3X1_616 ( .gnd(gnd), .vdd(vdd), .A(_3434_), .B(_2773_), .C(_2772_), .Y(_2778_) );
NAND3X1 NAND3X1_617 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_2778_), .C(_2777_), .Y(_2780_) );
NAND2X1 NAND2X1_344 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_237_), .B(_2780_), .Y(_2781_) );
AOI21X1 AOI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_2776_), .B(_2781_), .C(_2408_), .Y(_2782_) );
INVX1 INVX1_291 ( .gnd(gnd), .vdd(vdd), .A(_2408_), .Y(_2783_) );
NAND3X1 NAND3X1_618 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_237_), .B(_583_), .C(_2775_), .Y(_2784_) );
NAND2X1 NAND2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_2451_), .B(_2780_), .Y(_2785_) );
AOI21X1 AOI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_2784_), .B(_2785_), .C(_2783_), .Y(_2786_) );
OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_2782_), .B(_2786_), .C(_2450_), .Y(_2787_) );
OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_2423_), .B(_2430_), .C(_2416_), .Y(_2788_) );
NAND3X1 NAND3X1_619 ( .gnd(gnd), .vdd(vdd), .A(_2783_), .B(_2784_), .C(_2785_), .Y(_2789_) );
NAND3X1 NAND3X1_620 ( .gnd(gnd), .vdd(vdd), .A(_2408_), .B(_2776_), .C(_2781_), .Y(_2791_) );
NAND3X1 NAND3X1_621 ( .gnd(gnd), .vdd(vdd), .A(_2789_), .B(_2791_), .C(_2788_), .Y(_2792_) );
NAND3X1 NAND3X1_622 ( .gnd(gnd), .vdd(vdd), .A(_3631_), .B(_2787_), .C(_2792_), .Y(_2793_) );
AOI21X1 AOI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_2789_), .B(_2791_), .C(_2788_), .Y(_2794_) );
NOR3X1 NOR3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_2782_), .B(_2450_), .C(_2786_), .Y(_2795_) );
OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_2795_), .B(_2794_), .C(_3442_), .Y(_2796_) );
NAND2X1 NAND2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_2793_), .B(_2796_), .Y(_2797_) );
NAND3X1 NAND3X1_623 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_253_), .B(_591_), .C(_2797_), .Y(_2798_) );
INVX1 INVX1_292 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_253_), .Y(_2799_) );
OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_2795_), .B(_2794_), .C(_3631_), .Y(_2800_) );
NAND3X1 NAND3X1_624 ( .gnd(gnd), .vdd(vdd), .A(_3442_), .B(_2787_), .C(_2792_), .Y(_2802_) );
NAND3X1 NAND3X1_625 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_2802_), .C(_2800_), .Y(_2803_) );
NAND2X1 NAND2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_2799_), .B(_2803_), .Y(_2804_) );
NAND3X1 NAND3X1_626 ( .gnd(gnd), .vdd(vdd), .A(_2448_), .B(_2798_), .C(_2804_), .Y(_2805_) );
INVX1 INVX1_293 ( .gnd(gnd), .vdd(vdd), .A(_2448_), .Y(_2806_) );
NAND2X1 NAND2X1_348 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_253_), .B(_2803_), .Y(_2807_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_2803_), .B(module_0_W_253_), .Y(_2808_) );
NAND3X1 NAND3X1_627 ( .gnd(gnd), .vdd(vdd), .A(_2806_), .B(_2807_), .C(_2808_), .Y(_2809_) );
NAND2X1 NAND2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_2805_), .B(_2809_), .Y(_2810_) );
XNOR2X1 XNOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_2810_), .B(_2446_), .Y(module_0_H_21_) );
AOI21X1 AOI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2798_), .B(_2804_), .C(_2448_), .Y(_2812_) );
AOI21X1 AOI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2446_), .B(_2805_), .C(_2812_), .Y(_2813_) );
INVX1 INVX1_294 ( .gnd(gnd), .vdd(vdd), .A(_2813_), .Y(_2814_) );
INVX1 INVX1_295 ( .gnd(gnd), .vdd(vdd), .A(_2807_), .Y(_2815_) );
OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_2786_), .B(_2450_), .C(_2789_), .Y(_2816_) );
OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_2767_), .B(_2765_), .C(_2760_), .Y(_2817_) );
OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_2454_), .B(_2742_), .C(_2745_), .Y(_2818_) );
OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_2723_), .B(_2721_), .C(_2716_), .Y(_2819_) );
INVX1 INVX1_296 ( .gnd(gnd), .vdd(vdd), .A(_2819_), .Y(_2820_) );
INVX1 INVX1_297 ( .gnd(gnd), .vdd(vdd), .A(_2717_), .Y(_2821_) );
OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_2697_), .B(_2458_), .C(_2700_), .Y(_2823_) );
INVX1 INVX1_298 ( .gnd(gnd), .vdd(vdd), .A(_2823_), .Y(_2824_) );
INVX1 INVX1_299 ( .gnd(gnd), .vdd(vdd), .A(_2687_), .Y(_2825_) );
OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_2675_), .B(_2462_), .C(_2678_), .Y(_2826_) );
INVX1 INVX1_300 ( .gnd(gnd), .vdd(vdd), .A(_2826_), .Y(_2827_) );
INVX1 INVX1_301 ( .gnd(gnd), .vdd(vdd), .A(_2665_), .Y(_2828_) );
OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_2653_), .B(_2465_), .C(_2656_), .Y(_2829_) );
NAND2X1 NAND2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_2627_), .B(_2640_), .Y(_2830_) );
INVX1 INVX1_302 ( .gnd(gnd), .vdd(vdd), .A(_2830_), .Y(_2831_) );
NAND2X1 NAND2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_2612_), .B(_2615_), .Y(_2832_) );
NAND2X1 NAND2X1_352 ( .gnd(gnd), .vdd(vdd), .A(_2591_), .B(_2594_), .Y(_2834_) );
NAND2X1 NAND2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_2571_), .B(_2573_), .Y(_2835_) );
NAND2X1 NAND2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_2542_), .B(_2556_), .Y(_2836_) );
NAND2X1 NAND2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_2528_), .B(_2530_), .Y(_2837_) );
OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_2506_), .B(_2507_), .C(_2503_), .Y(_2838_) );
INVX1 INVX1_303 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_30_), .Y(_2839_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_12_), .B(module_0_W_13_), .Y(_2840_) );
XNOR2X1 XNOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_2840_), .B(module_0_W_14_), .Y(_2841_) );
XNOR2X1 XNOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_981_), .B(module_0_W_10_), .Y(_2842_) );
XNOR2X1 XNOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_2842_), .B(_2841_), .Y(_2843_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_2843_), .B(_2839_), .Y(_2845_) );
NAND2X1 NAND2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2839_), .B(_2843_), .Y(_2846_) );
NAND2X1 NAND2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_2846_), .B(_2845_), .Y(_2847_) );
XNOR2X1 XNOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_2847_), .B(_2499_), .Y(_2848_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_2848_), .B(_2838_), .Y(_2849_) );
XNOR2X1 XNOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .B(_1040_), .Y(_2850_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_2849_), .B(_2850_), .Y(_2851_) );
NAND2X1 NAND2X1_358 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf3_), .B(_2851_), .Y(_2852_) );
INVX1 INVX1_304 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf2_), .Y(_2853_) );
XNOR2X1 XNOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_2849_), .B(_2850_), .Y(_2854_) );
NAND2X1 NAND2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_2853_), .B(_2854_), .Y(_2856_) );
NAND3X1 NAND3X1_628 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .B(_2856_), .C(_2852_), .Y(_2857_) );
NAND2X1 NAND2X1_360 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf1_), .B(_2854_), .Y(_2858_) );
NAND2X1 NAND2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2853_), .B(_2851_), .Y(_2859_) );
NAND3X1 NAND3X1_629 ( .gnd(gnd), .vdd(vdd), .A(_2520_), .B(_2858_), .C(_2859_), .Y(_2860_) );
NAND3X1 NAND3X1_630 ( .gnd(gnd), .vdd(vdd), .A(_2837_), .B(_2857_), .C(_2860_), .Y(_2861_) );
AOI21X1 AOI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .B(_2860_), .C(_2837_), .Y(_2862_) );
INVX1 INVX1_305 ( .gnd(gnd), .vdd(vdd), .A(_2862_), .Y(_2863_) );
XNOR2X1 XNOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1075_), .B(_1026_), .Y(_2864_) );
NAND3X1 NAND3X1_631 ( .gnd(gnd), .vdd(vdd), .A(_2861_), .B(_2864_), .C(_2863_), .Y(_2865_) );
INVX1 INVX1_306 ( .gnd(gnd), .vdd(vdd), .A(_2861_), .Y(_2867_) );
INVX1 INVX1_307 ( .gnd(gnd), .vdd(vdd), .A(_2864_), .Y(_2868_) );
OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_2867_), .B(_2862_), .C(_2868_), .Y(_2869_) );
NAND3X1 NAND3X1_632 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf3_), .B(_2865_), .C(_2869_), .Y(_2870_) );
INVX1 INVX1_308 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf2_), .Y(_2871_) );
OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_2867_), .B(_2862_), .C(_2864_), .Y(_2872_) );
NAND3X1 NAND3X1_633 ( .gnd(gnd), .vdd(vdd), .A(_2861_), .B(_2868_), .C(_2863_), .Y(_2873_) );
NAND3X1 NAND3X1_634 ( .gnd(gnd), .vdd(vdd), .A(_2871_), .B(_2873_), .C(_2872_), .Y(_2874_) );
NAND3X1 NAND3X1_635 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .B(_2870_), .C(_2874_), .Y(_2875_) );
NAND3X1 NAND3X1_636 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf1_), .B(_2873_), .C(_2872_), .Y(_2876_) );
NAND3X1 NAND3X1_637 ( .gnd(gnd), .vdd(vdd), .A(_2871_), .B(_2865_), .C(_2869_), .Y(_2878_) );
NAND3X1 NAND3X1_638 ( .gnd(gnd), .vdd(vdd), .A(_2541_), .B(_2876_), .C(_2878_), .Y(_2879_) );
NAND3X1 NAND3X1_639 ( .gnd(gnd), .vdd(vdd), .A(_2836_), .B(_2875_), .C(_2879_), .Y(_2880_) );
INVX1 INVX1_309 ( .gnd(gnd), .vdd(vdd), .A(_2836_), .Y(_2881_) );
NAND3X1 NAND3X1_640 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .B(_2876_), .C(_2878_), .Y(_2882_) );
NAND3X1 NAND3X1_641 ( .gnd(gnd), .vdd(vdd), .A(_2541_), .B(_2870_), .C(_2874_), .Y(_2883_) );
NAND3X1 NAND3X1_642 ( .gnd(gnd), .vdd(vdd), .A(_2881_), .B(_2882_), .C(_2883_), .Y(_2884_) );
XNOR2X1 XNOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1113_), .B(_1063_), .Y(_2885_) );
NAND3X1 NAND3X1_643 ( .gnd(gnd), .vdd(vdd), .A(_2885_), .B(_2880_), .C(_2884_), .Y(_2886_) );
AOI21X1 AOI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_2882_), .B(_2883_), .C(_2881_), .Y(_2887_) );
AOI21X1 AOI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_2875_), .B(_2879_), .C(_2836_), .Y(_2889_) );
INVX1 INVX1_310 ( .gnd(gnd), .vdd(vdd), .A(_2885_), .Y(_2890_) );
OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_2887_), .B(_2889_), .C(_2890_), .Y(_2891_) );
NAND3X1 NAND3X1_644 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf4_), .B(_2886_), .C(_2891_), .Y(_2892_) );
INVX1 INVX1_311 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf3_), .Y(_2893_) );
OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_2887_), .B(_2889_), .C(_2885_), .Y(_2894_) );
NAND3X1 NAND3X1_645 ( .gnd(gnd), .vdd(vdd), .A(_2890_), .B(_2880_), .C(_2884_), .Y(_2895_) );
NAND3X1 NAND3X1_646 ( .gnd(gnd), .vdd(vdd), .A(_2893_), .B(_2895_), .C(_2894_), .Y(_2896_) );
NAND3X1 NAND3X1_647 ( .gnd(gnd), .vdd(vdd), .A(_2566_), .B(_2892_), .C(_2896_), .Y(_2897_) );
NAND3X1 NAND3X1_648 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf2_), .B(_2895_), .C(_2894_), .Y(_2898_) );
NAND3X1 NAND3X1_649 ( .gnd(gnd), .vdd(vdd), .A(_2893_), .B(_2886_), .C(_2891_), .Y(_2900_) );
NAND3X1 NAND3X1_650 ( .gnd(gnd), .vdd(vdd), .A(_2563_), .B(_2898_), .C(_2900_), .Y(_2901_) );
NAND3X1 NAND3X1_651 ( .gnd(gnd), .vdd(vdd), .A(_2835_), .B(_2897_), .C(_2901_), .Y(_2902_) );
INVX1 INVX1_312 ( .gnd(gnd), .vdd(vdd), .A(_2835_), .Y(_2903_) );
NAND3X1 NAND3X1_652 ( .gnd(gnd), .vdd(vdd), .A(_2566_), .B(_2898_), .C(_2900_), .Y(_2904_) );
NAND3X1 NAND3X1_653 ( .gnd(gnd), .vdd(vdd), .A(_2563_), .B(_2892_), .C(_2896_), .Y(_2905_) );
NAND3X1 NAND3X1_654 ( .gnd(gnd), .vdd(vdd), .A(_2903_), .B(_2904_), .C(_2905_), .Y(_2906_) );
XNOR2X1 XNOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1152_), .B(_3729_), .Y(_2907_) );
NAND3X1 NAND3X1_655 ( .gnd(gnd), .vdd(vdd), .A(_2907_), .B(_2902_), .C(_2906_), .Y(_2908_) );
AOI21X1 AOI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_2904_), .B(_2905_), .C(_2903_), .Y(_2909_) );
AOI21X1 AOI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2897_), .B(_2901_), .C(_2835_), .Y(_2911_) );
INVX1 INVX1_313 ( .gnd(gnd), .vdd(vdd), .A(_2907_), .Y(_2912_) );
OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_2909_), .B(_2911_), .C(_2912_), .Y(_2913_) );
NAND3X1 NAND3X1_656 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf3_), .B(_2908_), .C(_2913_), .Y(_2914_) );
INVX1 INVX1_314 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf2_), .Y(_2915_) );
OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_2909_), .B(_2911_), .C(_2907_), .Y(_2916_) );
NAND3X1 NAND3X1_657 ( .gnd(gnd), .vdd(vdd), .A(_2912_), .B(_2902_), .C(_2906_), .Y(_2917_) );
NAND3X1 NAND3X1_658 ( .gnd(gnd), .vdd(vdd), .A(_2915_), .B(_2917_), .C(_2916_), .Y(_2918_) );
NAND3X1 NAND3X1_659 ( .gnd(gnd), .vdd(vdd), .A(_2587_), .B(_2914_), .C(_2918_), .Y(_2919_) );
NAND3X1 NAND3X1_660 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf1_), .B(_2917_), .C(_2916_), .Y(_2920_) );
NAND3X1 NAND3X1_661 ( .gnd(gnd), .vdd(vdd), .A(_2915_), .B(_2908_), .C(_2913_), .Y(_2922_) );
NAND3X1 NAND3X1_662 ( .gnd(gnd), .vdd(vdd), .A(_2584_), .B(_2920_), .C(_2922_), .Y(_2923_) );
NAND3X1 NAND3X1_663 ( .gnd(gnd), .vdd(vdd), .A(_2834_), .B(_2919_), .C(_2923_), .Y(_2924_) );
INVX2 INVX2_70 ( .gnd(gnd), .vdd(vdd), .A(_2834_), .Y(_2925_) );
AOI21X1 AOI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_2920_), .B(_2922_), .C(_2584_), .Y(_2926_) );
AOI21X1 AOI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_2914_), .B(_2918_), .C(_2587_), .Y(_2927_) );
OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .B(_2927_), .C(_2925_), .Y(_2928_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1193_), .B(_1154_), .Y(_2929_) );
NAND3X1 NAND3X1_664 ( .gnd(gnd), .vdd(vdd), .A(_2924_), .B(_2929_), .C(_2928_), .Y(_2930_) );
NOR3X1 NOR3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .B(_2925_), .C(_2927_), .Y(_2931_) );
AOI21X1 AOI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_2919_), .B(_2923_), .C(_2834_), .Y(_2933_) );
INVX1 INVX1_315 ( .gnd(gnd), .vdd(vdd), .A(_2929_), .Y(_2934_) );
OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_2931_), .B(_2933_), .C(_2934_), .Y(_2935_) );
NAND3X1 NAND3X1_665 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf4_), .B(_2930_), .C(_2935_), .Y(_2936_) );
INVX1 INVX1_316 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf3_), .Y(_2937_) );
OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_2931_), .B(_2933_), .C(_2929_), .Y(_2938_) );
NAND3X1 NAND3X1_666 ( .gnd(gnd), .vdd(vdd), .A(_2924_), .B(_2934_), .C(_2928_), .Y(_2939_) );
NAND3X1 NAND3X1_667 ( .gnd(gnd), .vdd(vdd), .A(_2937_), .B(_2939_), .C(_2938_), .Y(_2940_) );
NAND3X1 NAND3X1_668 ( .gnd(gnd), .vdd(vdd), .A(_2608_), .B(_2936_), .C(_2940_), .Y(_2941_) );
NAND3X1 NAND3X1_669 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf2_), .B(_2939_), .C(_2938_), .Y(_2942_) );
NAND3X1 NAND3X1_670 ( .gnd(gnd), .vdd(vdd), .A(_2937_), .B(_2930_), .C(_2935_), .Y(_2944_) );
NAND3X1 NAND3X1_671 ( .gnd(gnd), .vdd(vdd), .A(_2605_), .B(_2942_), .C(_2944_), .Y(_2945_) );
NAND3X1 NAND3X1_672 ( .gnd(gnd), .vdd(vdd), .A(_2832_), .B(_2941_), .C(_2945_), .Y(_2946_) );
INVX1 INVX1_317 ( .gnd(gnd), .vdd(vdd), .A(_2832_), .Y(_2947_) );
NAND3X1 NAND3X1_673 ( .gnd(gnd), .vdd(vdd), .A(_2608_), .B(_2942_), .C(_2944_), .Y(_2948_) );
NAND3X1 NAND3X1_674 ( .gnd(gnd), .vdd(vdd), .A(_2605_), .B(_2936_), .C(_2940_), .Y(_2949_) );
NAND3X1 NAND3X1_675 ( .gnd(gnd), .vdd(vdd), .A(_2947_), .B(_2948_), .C(_2949_), .Y(_2950_) );
XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1233_), .B(_1195_), .Y(_2951_) );
INVX1 INVX1_318 ( .gnd(gnd), .vdd(vdd), .A(_2951_), .Y(_2952_) );
NAND3X1 NAND3X1_676 ( .gnd(gnd), .vdd(vdd), .A(_2952_), .B(_2946_), .C(_2950_), .Y(_2953_) );
AOI21X1 AOI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_2948_), .B(_2949_), .C(_2947_), .Y(_2955_) );
AOI21X1 AOI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_2941_), .B(_2945_), .C(_2832_), .Y(_2956_) );
OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_2955_), .B(_2956_), .C(_2951_), .Y(_2957_) );
NAND3X1 NAND3X1_677 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf3_), .B(_2953_), .C(_2957_), .Y(_2958_) );
INVX1 INVX1_319 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf2_), .Y(_2959_) );
NAND3X1 NAND3X1_678 ( .gnd(gnd), .vdd(vdd), .A(_2951_), .B(_2946_), .C(_2950_), .Y(_2960_) );
OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_2955_), .B(_2956_), .C(_2952_), .Y(_2961_) );
NAND3X1 NAND3X1_679 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .B(_2960_), .C(_2961_), .Y(_2962_) );
NAND3X1 NAND3X1_680 ( .gnd(gnd), .vdd(vdd), .A(_2630_), .B(_2958_), .C(_2962_), .Y(_2963_) );
NAND3X1 NAND3X1_681 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf1_), .B(_2960_), .C(_2961_), .Y(_2964_) );
NAND3X1 NAND3X1_682 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .B(_2953_), .C(_2957_), .Y(_2966_) );
NAND3X1 NAND3X1_683 ( .gnd(gnd), .vdd(vdd), .A(_2626_), .B(_2964_), .C(_2966_), .Y(_2967_) );
AOI21X1 AOI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_2963_), .B(_2967_), .C(_2831_), .Y(_2968_) );
NAND3X1 NAND3X1_684 ( .gnd(gnd), .vdd(vdd), .A(_2630_), .B(_2964_), .C(_2966_), .Y(_2969_) );
NAND3X1 NAND3X1_685 ( .gnd(gnd), .vdd(vdd), .A(_2626_), .B(_2958_), .C(_2962_), .Y(_2970_) );
AOI21X1 AOI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_2969_), .B(_2970_), .C(_2830_), .Y(_2971_) );
OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_2968_), .B(_2971_), .C(_1235_), .Y(_2972_) );
INVX1 INVX1_320 ( .gnd(gnd), .vdd(vdd), .A(_1235_), .Y(_2973_) );
NAND3X1 NAND3X1_686 ( .gnd(gnd), .vdd(vdd), .A(_2830_), .B(_2969_), .C(_2970_), .Y(_2974_) );
NAND3X1 NAND3X1_687 ( .gnd(gnd), .vdd(vdd), .A(_2963_), .B(_2967_), .C(_2831_), .Y(_2975_) );
NAND3X1 NAND3X1_688 ( .gnd(gnd), .vdd(vdd), .A(_2973_), .B(_2974_), .C(_2975_), .Y(_2977_) );
NAND3X1 NAND3X1_689 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .B(_2977_), .C(_2972_), .Y(_2978_) );
NAND2X1 NAND2X1_362 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_142_), .B(_2978_), .Y(_2979_) );
INVX1 INVX1_321 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_142_), .Y(_2980_) );
OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_2968_), .B(_2971_), .C(_2973_), .Y(_2981_) );
NAND3X1 NAND3X1_690 ( .gnd(gnd), .vdd(vdd), .A(_1235_), .B(_2974_), .C(_2975_), .Y(_2982_) );
NAND2X1 NAND2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2981_), .Y(_2983_) );
NAND3X1 NAND3X1_691 ( .gnd(gnd), .vdd(vdd), .A(_2980_), .B(_1274_), .C(_2983_), .Y(_2984_) );
NAND3X1 NAND3X1_692 ( .gnd(gnd), .vdd(vdd), .A(_2643_), .B(_2984_), .C(_2979_), .Y(_2985_) );
INVX1 INVX1_322 ( .gnd(gnd), .vdd(vdd), .A(_2643_), .Y(_2986_) );
NAND3X1 NAND3X1_693 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_142_), .B(_1274_), .C(_2983_), .Y(_2988_) );
NAND2X1 NAND2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_2980_), .B(_2978_), .Y(_2989_) );
NAND3X1 NAND3X1_694 ( .gnd(gnd), .vdd(vdd), .A(_2986_), .B(_2988_), .C(_2989_), .Y(_2990_) );
NAND3X1 NAND3X1_695 ( .gnd(gnd), .vdd(vdd), .A(_2829_), .B(_2985_), .C(_2990_), .Y(_2991_) );
INVX1 INVX1_323 ( .gnd(gnd), .vdd(vdd), .A(_2829_), .Y(_2992_) );
NAND3X1 NAND3X1_696 ( .gnd(gnd), .vdd(vdd), .A(_2986_), .B(_2984_), .C(_2979_), .Y(_2993_) );
NAND3X1 NAND3X1_697 ( .gnd(gnd), .vdd(vdd), .A(_2643_), .B(_2988_), .C(_2989_), .Y(_2994_) );
NAND3X1 NAND3X1_698 ( .gnd(gnd), .vdd(vdd), .A(_2992_), .B(_2993_), .C(_2994_), .Y(_2995_) );
NAND3X1 NAND3X1_699 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_2991_), .C(_2995_), .Y(_2996_) );
AOI21X1 AOI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_2993_), .B(_2994_), .C(_2992_), .Y(_2997_) );
AOI21X1 AOI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_2985_), .B(_2990_), .C(_2829_), .Y(_2999_) );
OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2997_), .B(_2999_), .C(_961_), .Y(_3000_) );
NAND3X1 NAND3X1_700 ( .gnd(gnd), .vdd(vdd), .A(_1308_), .B(_2996_), .C(_3000_), .Y(_3001_) );
NAND2X1 NAND2X1_365 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_158_), .B(_3001_), .Y(_3002_) );
INVX1 INVX1_324 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_158_), .Y(_3003_) );
NAND2X1 NAND2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_2991_), .B(_2995_), .Y(_3004_) );
AOI21X1 AOI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_961_), .B(_3004_), .C(_1309_), .Y(_3005_) );
NAND3X1 NAND3X1_701 ( .gnd(gnd), .vdd(vdd), .A(_3003_), .B(_2996_), .C(_3005_), .Y(_3006_) );
NAND3X1 NAND3X1_702 ( .gnd(gnd), .vdd(vdd), .A(_2828_), .B(_3006_), .C(_3002_), .Y(_3007_) );
NAND3X1 NAND3X1_703 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_158_), .B(_2996_), .C(_3005_), .Y(_3008_) );
NAND2X1 NAND2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_3003_), .B(_3001_), .Y(_3010_) );
NAND3X1 NAND3X1_704 ( .gnd(gnd), .vdd(vdd), .A(_2665_), .B(_3008_), .C(_3010_), .Y(_3011_) );
AOI21X1 AOI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_3007_), .B(_3011_), .C(_2827_), .Y(_3012_) );
NAND3X1 NAND3X1_705 ( .gnd(gnd), .vdd(vdd), .A(_2665_), .B(_3006_), .C(_3002_), .Y(_3013_) );
NAND3X1 NAND3X1_706 ( .gnd(gnd), .vdd(vdd), .A(_2828_), .B(_3008_), .C(_3010_), .Y(_3014_) );
AOI21X1 AOI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_3013_), .B(_3014_), .C(_2826_), .Y(_3015_) );
OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_3012_), .B(_3015_), .C(_3574_), .Y(_3016_) );
NAND3X1 NAND3X1_707 ( .gnd(gnd), .vdd(vdd), .A(_2826_), .B(_3013_), .C(_3014_), .Y(_3017_) );
NAND3X1 NAND3X1_708 ( .gnd(gnd), .vdd(vdd), .A(_2827_), .B(_3007_), .C(_3011_), .Y(_3018_) );
NAND3X1 NAND3X1_709 ( .gnd(gnd), .vdd(vdd), .A(_3787_), .B(_3017_), .C(_3018_), .Y(_3019_) );
NAND3X1 NAND3X1_710 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_3019_), .C(_3016_), .Y(_3021_) );
NAND2X1 NAND2X1_368 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_174_), .B(_3021_), .Y(_3022_) );
INVX1 INVX1_325 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_174_), .Y(_3023_) );
OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_3012_), .B(_3015_), .C(_3787_), .Y(_3024_) );
NAND3X1 NAND3X1_711 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .B(_3017_), .C(_3018_), .Y(_3025_) );
NAND2X1 NAND2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_3025_), .B(_3024_), .Y(_3026_) );
NAND3X1 NAND3X1_712 ( .gnd(gnd), .vdd(vdd), .A(_3023_), .B(_1343_), .C(_3026_), .Y(_3027_) );
NAND3X1 NAND3X1_713 ( .gnd(gnd), .vdd(vdd), .A(_2825_), .B(_3027_), .C(_3022_), .Y(_3028_) );
NAND3X1 NAND3X1_714 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_174_), .B(_1343_), .C(_3026_), .Y(_3029_) );
NAND2X1 NAND2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_3023_), .B(_3021_), .Y(_3030_) );
NAND3X1 NAND3X1_715 ( .gnd(gnd), .vdd(vdd), .A(_2687_), .B(_3029_), .C(_3030_), .Y(_3032_) );
AOI21X1 AOI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_3028_), .B(_3032_), .C(_2824_), .Y(_3033_) );
NAND3X1 NAND3X1_716 ( .gnd(gnd), .vdd(vdd), .A(_2687_), .B(_3027_), .C(_3022_), .Y(_3034_) );
NAND3X1 NAND3X1_717 ( .gnd(gnd), .vdd(vdd), .A(_2825_), .B(_3029_), .C(_3030_), .Y(_3035_) );
AOI21X1 AOI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_3034_), .B(_3035_), .C(_2823_), .Y(_3036_) );
OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_3036_), .B(_3033_), .C(_3584_), .Y(_3037_) );
NAND3X1 NAND3X1_718 ( .gnd(gnd), .vdd(vdd), .A(_2823_), .B(_3034_), .C(_3035_), .Y(_3038_) );
NAND3X1 NAND3X1_719 ( .gnd(gnd), .vdd(vdd), .A(_3028_), .B(_2824_), .C(_3032_), .Y(_3039_) );
NAND3X1 NAND3X1_720 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_3038_), .C(_3039_), .Y(_3040_) );
NAND3X1 NAND3X1_721 ( .gnd(gnd), .vdd(vdd), .A(_1381_), .B(_3040_), .C(_3037_), .Y(_3041_) );
NAND2X1 NAND2X1_371 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_190_), .B(_3041_), .Y(_3043_) );
INVX1 INVX1_326 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_190_), .Y(_3044_) );
OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_3036_), .B(_3033_), .C(_956_), .Y(_3045_) );
NAND3X1 NAND3X1_722 ( .gnd(gnd), .vdd(vdd), .A(_3584_), .B(_3038_), .C(_3039_), .Y(_3046_) );
NAND2X1 NAND2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_3046_), .B(_3045_), .Y(_3047_) );
NAND3X1 NAND3X1_723 ( .gnd(gnd), .vdd(vdd), .A(_3044_), .B(_1381_), .C(_3047_), .Y(_3048_) );
NAND3X1 NAND3X1_724 ( .gnd(gnd), .vdd(vdd), .A(_2821_), .B(_3048_), .C(_3043_), .Y(_3049_) );
NAND3X1 NAND3X1_725 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_190_), .B(_1381_), .C(_3047_), .Y(_3050_) );
NAND2X1 NAND2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_3044_), .B(_3041_), .Y(_3051_) );
NAND3X1 NAND3X1_726 ( .gnd(gnd), .vdd(vdd), .A(_2717_), .B(_3050_), .C(_3051_), .Y(_3052_) );
AOI21X1 AOI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_3049_), .B(_3052_), .C(_2820_), .Y(_3054_) );
NAND3X1 NAND3X1_727 ( .gnd(gnd), .vdd(vdd), .A(_2717_), .B(_3048_), .C(_3043_), .Y(_3055_) );
NAND3X1 NAND3X1_728 ( .gnd(gnd), .vdd(vdd), .A(_2821_), .B(_3050_), .C(_3051_), .Y(_3056_) );
AOI21X1 AOI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .B(_3056_), .C(_2819_), .Y(_3057_) );
OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_3054_), .B(_3057_), .C(_952_), .Y(_3058_) );
NAND3X1 NAND3X1_729 ( .gnd(gnd), .vdd(vdd), .A(_2819_), .B(_3055_), .C(_3056_), .Y(_3059_) );
NAND3X1 NAND3X1_730 ( .gnd(gnd), .vdd(vdd), .A(_3049_), .B(_3052_), .C(_2820_), .Y(_3060_) );
NAND3X1 NAND3X1_731 ( .gnd(gnd), .vdd(vdd), .A(_953_), .B(_3059_), .C(_3060_), .Y(_3061_) );
NAND3X1 NAND3X1_732 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .B(_3061_), .C(_3058_), .Y(_3062_) );
NAND2X1 NAND2X1_374 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_206_), .B(_3062_), .Y(_3063_) );
INVX1 INVX1_327 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_206_), .Y(_3065_) );
NAND3X1 NAND3X1_733 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_3059_), .C(_3060_), .Y(_3066_) );
OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_3054_), .B(_3057_), .C(_953_), .Y(_3067_) );
NAND2X1 NAND2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_3066_), .B(_3067_), .Y(_3068_) );
NAND3X1 NAND3X1_734 ( .gnd(gnd), .vdd(vdd), .A(_3065_), .B(_1417_), .C(_3068_), .Y(_3069_) );
NAND3X1 NAND3X1_735 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .B(_3069_), .C(_3063_), .Y(_3070_) );
INVX1 INVX1_328 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .Y(_3071_) );
NAND3X1 NAND3X1_736 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_206_), .B(_1417_), .C(_3068_), .Y(_3072_) );
NAND2X1 NAND2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_3065_), .B(_3062_), .Y(_3073_) );
NAND3X1 NAND3X1_737 ( .gnd(gnd), .vdd(vdd), .A(_3071_), .B(_3072_), .C(_3073_), .Y(_3074_) );
NAND3X1 NAND3X1_738 ( .gnd(gnd), .vdd(vdd), .A(_2818_), .B(_3070_), .C(_3074_), .Y(_3076_) );
AOI21X1 AOI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_2747_), .B(_2744_), .C(_2738_), .Y(_3077_) );
AOI21X1 AOI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_3072_), .B(_3073_), .C(_3071_), .Y(_3078_) );
AOI21X1 AOI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_3069_), .B(_3063_), .C(_2732_), .Y(_3079_) );
OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_3078_), .B(_3079_), .C(_3077_), .Y(_3080_) );
NAND3X1 NAND3X1_739 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(_3076_), .C(_3080_), .Y(_3081_) );
NOR3X1 NOR3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_3078_), .B(_3077_), .C(_3079_), .Y(_3082_) );
AOI21X1 AOI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_3070_), .B(_3074_), .C(_2818_), .Y(_3083_) );
OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_3082_), .B(_3083_), .C(_3602_), .Y(_3084_) );
NAND3X1 NAND3X1_740 ( .gnd(gnd), .vdd(vdd), .A(_1454_), .B(_3081_), .C(_3084_), .Y(_3085_) );
NAND2X1 NAND2X1_377 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_222_), .B(_3085_), .Y(_3087_) );
INVX1 INVX1_329 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_222_), .Y(_3088_) );
NAND2X1 NAND2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_3076_), .B(_3080_), .Y(_3089_) );
AOI21X1 AOI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_3602_), .B(_3089_), .C(_1455_), .Y(_3090_) );
NAND3X1 NAND3X1_741 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_3081_), .C(_3090_), .Y(_3091_) );
NAND3X1 NAND3X1_742 ( .gnd(gnd), .vdd(vdd), .A(_2761_), .B(_3091_), .C(_3087_), .Y(_3092_) );
INVX1 INVX1_330 ( .gnd(gnd), .vdd(vdd), .A(_2761_), .Y(_3093_) );
NAND3X1 NAND3X1_743 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_222_), .B(_3081_), .C(_3090_), .Y(_3094_) );
NAND2X1 NAND2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_3085_), .Y(_3095_) );
NAND3X1 NAND3X1_744 ( .gnd(gnd), .vdd(vdd), .A(_3093_), .B(_3094_), .C(_3095_), .Y(_3096_) );
NAND3X1 NAND3X1_745 ( .gnd(gnd), .vdd(vdd), .A(_2817_), .B(_3092_), .C(_3096_), .Y(_3098_) );
AOI21X1 AOI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_2763_), .B(_2452_), .C(_2766_), .Y(_3099_) );
NAND3X1 NAND3X1_746 ( .gnd(gnd), .vdd(vdd), .A(_3093_), .B(_3091_), .C(_3087_), .Y(_3100_) );
NAND3X1 NAND3X1_747 ( .gnd(gnd), .vdd(vdd), .A(_2761_), .B(_3094_), .C(_3095_), .Y(_3101_) );
NAND3X1 NAND3X1_748 ( .gnd(gnd), .vdd(vdd), .A(_3099_), .B(_3100_), .C(_3101_), .Y(_3102_) );
NAND3X1 NAND3X1_749 ( .gnd(gnd), .vdd(vdd), .A(_946_), .B(_3098_), .C(_3102_), .Y(_3103_) );
AOI21X1 AOI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_3100_), .B(_3101_), .C(_3099_), .Y(_3104_) );
AOI21X1 AOI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3096_), .C(_2817_), .Y(_3105_) );
OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_3104_), .B(_3105_), .C(_945_), .Y(_3106_) );
NAND3X1 NAND3X1_750 ( .gnd(gnd), .vdd(vdd), .A(_1491_), .B(_3103_), .C(_3106_), .Y(_3107_) );
NAND2X1 NAND2X1_380 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_238_), .B(_3107_), .Y(_3109_) );
INVX1 INVX1_331 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_238_), .Y(_3110_) );
NAND2X1 NAND2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_3098_), .B(_3102_), .Y(_3111_) );
AOI21X1 AOI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_945_), .B(_3111_), .C(_1492_), .Y(_3112_) );
NAND3X1 NAND3X1_751 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .B(_3103_), .C(_3112_), .Y(_3113_) );
NAND3X1 NAND3X1_752 ( .gnd(gnd), .vdd(vdd), .A(_2776_), .B(_3113_), .C(_3109_), .Y(_3114_) );
INVX2 INVX2_71 ( .gnd(gnd), .vdd(vdd), .A(_2776_), .Y(_3115_) );
NAND3X1 NAND3X1_753 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_238_), .B(_3103_), .C(_3112_), .Y(_3116_) );
NAND2X1 NAND2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .B(_3107_), .Y(_3117_) );
NAND3X1 NAND3X1_754 ( .gnd(gnd), .vdd(vdd), .A(_3115_), .B(_3116_), .C(_3117_), .Y(_3118_) );
NAND3X1 NAND3X1_755 ( .gnd(gnd), .vdd(vdd), .A(_3114_), .B(_3118_), .C(_2816_), .Y(_3120_) );
AOI21X1 AOI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_2791_), .B(_2788_), .C(_2782_), .Y(_3121_) );
AOI21X1 AOI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_3116_), .B(_3117_), .C(_3115_), .Y(_3122_) );
AOI21X1 AOI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .B(_3109_), .C(_2776_), .Y(_3123_) );
OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_3122_), .B(_3123_), .C(_3121_), .Y(_3124_) );
NAND3X1 NAND3X1_756 ( .gnd(gnd), .vdd(vdd), .A(_3852_), .B(_3120_), .C(_3124_), .Y(_3125_) );
NAND3X1 NAND3X1_757 ( .gnd(gnd), .vdd(vdd), .A(_3115_), .B(_3113_), .C(_3109_), .Y(_3126_) );
NAND3X1 NAND3X1_758 ( .gnd(gnd), .vdd(vdd), .A(_2776_), .B(_3116_), .C(_3117_), .Y(_3127_) );
AOI21X1 AOI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_3126_), .B(_3127_), .C(_3121_), .Y(_3128_) );
AOI21X1 AOI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_3114_), .B(_3118_), .C(_2816_), .Y(_3129_) );
OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_3128_), .B(_3129_), .C(_3624_), .Y(_3131_) );
NAND3X1 NAND3X1_759 ( .gnd(gnd), .vdd(vdd), .A(_1526_), .B(_3125_), .C(_3131_), .Y(_3132_) );
NAND2X1 NAND2X1_383 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_254_), .B(_3132_), .Y(_3133_) );
INVX1 INVX1_332 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_254_), .Y(_3134_) );
NAND2X1 NAND2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_3120_), .B(_3124_), .Y(_3135_) );
AOI21X1 AOI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_3624_), .B(_3135_), .C(_1527_), .Y(_3136_) );
NAND3X1 NAND3X1_760 ( .gnd(gnd), .vdd(vdd), .A(_3134_), .B(_3125_), .C(_3136_), .Y(_3137_) );
NAND3X1 NAND3X1_761 ( .gnd(gnd), .vdd(vdd), .A(_2815_), .B(_3137_), .C(_3133_), .Y(_3138_) );
INVX1 INVX1_333 ( .gnd(gnd), .vdd(vdd), .A(_3138_), .Y(_3139_) );
AOI21X1 AOI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_3137_), .B(_3133_), .C(_2815_), .Y(_3140_) );
OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_3139_), .B(_3140_), .C(_2814_), .Y(_3142_) );
INVX1 INVX1_334 ( .gnd(gnd), .vdd(vdd), .A(_3140_), .Y(_3143_) );
NAND3X1 NAND3X1_762 ( .gnd(gnd), .vdd(vdd), .A(_2813_), .B(_3138_), .C(_3143_), .Y(_3144_) );
NAND2X1 NAND2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_3142_), .B(_3144_), .Y(module_0_H_22_) );
OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_2813_), .B(_3140_), .C(_3138_), .Y(_3145_) );
AOI21X1 AOI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_3125_), .B(_3136_), .C(_3134_), .Y(_3146_) );
INVX1 INVX1_335 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_255_), .Y(_3147_) );
OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_3121_), .B(_3123_), .C(_3114_), .Y(_3148_) );
INVX1 INVX1_336 ( .gnd(gnd), .vdd(vdd), .A(_3148_), .Y(_3149_) );
NAND2X1 NAND2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3098_), .Y(_3150_) );
OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_3079_), .B(_3077_), .C(_3070_), .Y(_3152_) );
NAND2X1 NAND2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .B(_3059_), .Y(_3153_) );
NAND2X1 NAND2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_3034_), .B(_3038_), .Y(_3154_) );
INVX1 INVX1_337 ( .gnd(gnd), .vdd(vdd), .A(_3154_), .Y(_3155_) );
NAND2X1 NAND2X1_389 ( .gnd(gnd), .vdd(vdd), .A(_3013_), .B(_3017_), .Y(_3156_) );
NAND2X1 NAND2X1_390 ( .gnd(gnd), .vdd(vdd), .A(_2985_), .B(_2991_), .Y(_3157_) );
NAND2X1 NAND2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_2969_), .B(_2974_), .Y(_3158_) );
INVX1 INVX1_338 ( .gnd(gnd), .vdd(vdd), .A(_3158_), .Y(_3159_) );
INVX1 INVX1_339 ( .gnd(gnd), .vdd(vdd), .A(_2964_), .Y(_3160_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_3758_), .B(_3760_), .Y(_3161_) );
NAND2X1 NAND2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_2941_), .B(_2946_), .Y(_3163_) );
INVX1 INVX1_340 ( .gnd(gnd), .vdd(vdd), .A(_3163_), .Y(_3164_) );
OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_2927_), .B(_2925_), .C(_2919_), .Y(_3165_) );
INVX1 INVX1_341 ( .gnd(gnd), .vdd(vdd), .A(_3740_), .Y(_3166_) );
NAND2X1 NAND2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_2897_), .B(_2902_), .Y(_3167_) );
INVX1 INVX1_342 ( .gnd(gnd), .vdd(vdd), .A(_3167_), .Y(_3168_) );
NAND2X1 NAND2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_2875_), .B(_2880_), .Y(_3169_) );
INVX1 INVX1_343 ( .gnd(gnd), .vdd(vdd), .A(_1778_), .Y(_3170_) );
XNOR2X1 XNOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_2870_), .B(_3170_), .Y(_3171_) );
INVX1 INVX1_344 ( .gnd(gnd), .vdd(vdd), .A(_3171_), .Y(_3172_) );
INVX1 INVX1_345 ( .gnd(gnd), .vdd(vdd), .A(_2837_), .Y(_3174_) );
NAND2X1 NAND2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .B(_2860_), .Y(_3175_) );
OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_3175_), .B(_3174_), .C(_2857_), .Y(_3176_) );
INVX1 INVX1_346 ( .gnd(gnd), .vdd(vdd), .A(_3176_), .Y(_3177_) );
INVX1 INVX1_347 ( .gnd(gnd), .vdd(vdd), .A(_2852_), .Y(_3178_) );
OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_2508_), .B(_2513_), .C(_2848_), .Y(_3179_) );
OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_2502_), .B(_2847_), .C(_3179_), .Y(_3180_) );
INVX1 INVX1_348 ( .gnd(gnd), .vdd(vdd), .A(_3180_), .Y(_3181_) );
OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_12_), .B(module_0_W_13_), .C(module_0_W_14_), .Y(_3182_) );
XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_11_), .B(module_0_W_15_), .Y(_3183_) );
XNOR2X1 XNOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_3183_), .B(_3182_), .Y(_3185_) );
XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .B(module_0_W_31_), .Y(_3186_) );
XNOR2X1 XNOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_3186_), .B(_3185_), .Y(_3187_) );
XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_2845_), .B(_3187_), .Y(_3188_) );
XNOR2X1 XNOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_3188_), .B(_1574_), .Y(_3189_) );
XNOR2X1 XNOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1742_), .B(bloque_datos[15]), .Y(_3190_) );
XNOR2X1 XNOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_3189_), .B(_3190_), .Y(_3191_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_3181_), .B(_3191_), .Y(_3192_) );
NAND2X1 NAND2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_3181_), .B(_3191_), .Y(_3193_) );
INVX1 INVX1_349 ( .gnd(gnd), .vdd(vdd), .A(_3193_), .Y(_3194_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_3194_), .B(_3192_), .Y(_3196_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_3178_), .B(_3196_), .Y(_3197_) );
INVX1 INVX1_350 ( .gnd(gnd), .vdd(vdd), .A(_3197_), .Y(_3198_) );
OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_3194_), .B(_3192_), .C(_3178_), .Y(_3199_) );
XNOR2X1 XNOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1756_), .B(_1580_), .Y(_3200_) );
INVX1 INVX1_351 ( .gnd(gnd), .vdd(vdd), .A(_3200_), .Y(_3201_) );
NAND3X1 NAND3X1_763 ( .gnd(gnd), .vdd(vdd), .A(_3199_), .B(_3201_), .C(_3198_), .Y(_3202_) );
AOI21X1 AOI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_3199_), .B(_3198_), .C(_3201_), .Y(_3203_) );
INVX1 INVX1_352 ( .gnd(gnd), .vdd(vdd), .A(_3203_), .Y(_3204_) );
NAND2X1 NAND2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_3202_), .B(_3204_), .Y(_3205_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf3_), .B(_3205_), .Y(_3207_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_3205_), .B(bloque_datos_31_bF_buf2_), .Y(_3208_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_3207_), .B(_3208_), .Y(_3209_) );
NAND2X1 NAND2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_3177_), .B(_3209_), .Y(_3210_) );
OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_3208_), .B(_3207_), .C(_3176_), .Y(_3211_) );
XOR2X1 XOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1595_), .B(bloque_datos_47_bF_buf3_), .Y(_3212_) );
NAND3X1 NAND3X1_764 ( .gnd(gnd), .vdd(vdd), .A(_3211_), .B(_3212_), .C(_3210_), .Y(_3213_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_3209_), .B(_3177_), .Y(_3214_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_3177_), .B(_3209_), .Y(_3215_) );
INVX1 INVX1_353 ( .gnd(gnd), .vdd(vdd), .A(_3212_), .Y(_3216_) );
OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_3214_), .B(_3215_), .C(_3216_), .Y(_3218_) );
AOI21X1 AOI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_3218_), .C(_3172_), .Y(_3219_) );
INVX1 INVX1_354 ( .gnd(gnd), .vdd(vdd), .A(_3219_), .Y(_3220_) );
NAND3X1 NAND3X1_765 ( .gnd(gnd), .vdd(vdd), .A(_3172_), .B(_3213_), .C(_3218_), .Y(_3221_) );
NAND3X1 NAND3X1_766 ( .gnd(gnd), .vdd(vdd), .A(_3169_), .B(_3221_), .C(_3220_), .Y(_3222_) );
INVX1 INVX1_355 ( .gnd(gnd), .vdd(vdd), .A(_3169_), .Y(_3223_) );
INVX1 INVX1_356 ( .gnd(gnd), .vdd(vdd), .A(_3221_), .Y(_3224_) );
OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_3224_), .B(_3219_), .C(_3223_), .Y(_3225_) );
OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .B(_1603_), .C(_3896_), .Y(_3226_) );
NAND2X1 NAND2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_3725_), .B(_1730_), .Y(_3227_) );
NAND2X1 NAND2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_3227_), .Y(_3229_) );
AOI21X1 AOI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_3225_), .B(_3222_), .C(_3229_), .Y(_3230_) );
NAND3X1 NAND3X1_767 ( .gnd(gnd), .vdd(vdd), .A(_3223_), .B(_3221_), .C(_3220_), .Y(_3231_) );
OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_3224_), .B(_3219_), .C(_3169_), .Y(_3232_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_3227_), .C(_3231_), .D(_3232_), .Y(_3233_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_3230_), .B(_3233_), .Y(_3234_) );
XNOR2X1 XNOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_2892_), .B(bloque_datos[63]), .Y(_3235_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_3234_), .B(_3235_), .Y(_3236_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_3235_), .B(_3234_), .Y(_3237_) );
OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_3236_), .B(_3237_), .C(_3168_), .Y(_3238_) );
NAND2X1 NAND2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_3235_), .B(_3234_), .Y(_3240_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_3234_), .B(_3235_), .Y(_3241_) );
NAND3X1 NAND3X1_768 ( .gnd(gnd), .vdd(vdd), .A(_3167_), .B(_3240_), .C(_3241_), .Y(_3242_) );
NAND3X1 NAND3X1_769 ( .gnd(gnd), .vdd(vdd), .A(_3166_), .B(_3238_), .C(_3242_), .Y(_3243_) );
NAND3X1 NAND3X1_770 ( .gnd(gnd), .vdd(vdd), .A(_3168_), .B(_3240_), .C(_3241_), .Y(_3244_) );
OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_3236_), .B(_3237_), .C(_3167_), .Y(_3245_) );
NAND3X1 NAND3X1_771 ( .gnd(gnd), .vdd(vdd), .A(_3740_), .B(_3245_), .C(_3244_), .Y(_3246_) );
NAND2X1 NAND2X1_402 ( .gnd(gnd), .vdd(vdd), .A(_3243_), .B(_3246_), .Y(_3247_) );
XOR2X1 XOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1728_), .B(bloque_datos_79_bF_buf3_), .Y(_3248_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_2914_), .B(_3248_), .Y(_3249_) );
INVX1 INVX1_357 ( .gnd(gnd), .vdd(vdd), .A(_3249_), .Y(_3251_) );
NAND2X1 NAND2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_2914_), .B(_3248_), .Y(_3252_) );
NAND2X1 NAND2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_3252_), .B(_3251_), .Y(_3253_) );
NAND2X1 NAND2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_3253_), .B(_3247_), .Y(_3254_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_3247_), .B(_3253_), .Y(_3255_) );
NAND3X1 NAND3X1_772 ( .gnd(gnd), .vdd(vdd), .A(_3165_), .B(_3254_), .C(_3255_), .Y(_3256_) );
INVX1 INVX1_358 ( .gnd(gnd), .vdd(vdd), .A(_3165_), .Y(_3257_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_3247_), .B(_3253_), .Y(_3258_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_3253_), .B(_3247_), .Y(_3259_) );
OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_3258_), .B(_3259_), .C(_3257_), .Y(_3260_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_3746_), .B(_3748_), .Y(_3262_) );
XNOR2X1 XNOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1726_), .B(_3262_), .Y(_3263_) );
INVX1 INVX1_359 ( .gnd(gnd), .vdd(vdd), .A(_3263_), .Y(_3264_) );
AOI21X1 AOI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_3260_), .B(_3256_), .C(_3264_), .Y(_3265_) );
NAND3X1 NAND3X1_773 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_3254_), .C(_3255_), .Y(_3266_) );
OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_3258_), .B(_3259_), .C(_3165_), .Y(_3267_) );
AOI21X1 AOI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_3267_), .B(_3266_), .C(_3263_), .Y(_3268_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_3265_), .B(_3268_), .Y(_3269_) );
NAND2X1 NAND2X1_406 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf3_), .B(_2936_), .Y(_3270_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf2_), .B(_2936_), .Y(_3271_) );
INVX1 INVX1_360 ( .gnd(gnd), .vdd(vdd), .A(_3271_), .Y(_3273_) );
NAND2X1 NAND2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_3270_), .B(_3273_), .Y(_3274_) );
NAND2X1 NAND2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_3274_), .B(_3269_), .Y(_3275_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_3269_), .B(_3274_), .Y(_3276_) );
NAND3X1 NAND3X1_774 ( .gnd(gnd), .vdd(vdd), .A(_3164_), .B(_3275_), .C(_3276_), .Y(_3277_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_3269_), .B(_3274_), .Y(_3278_) );
NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_3274_), .B(_3269_), .Y(_3279_) );
OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_3278_), .B(_3279_), .C(_3163_), .Y(_3280_) );
AOI21X1 AOI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_3280_), .B(_3277_), .C(_3161_), .Y(_3281_) );
INVX1 INVX1_361 ( .gnd(gnd), .vdd(vdd), .A(_3161_), .Y(_3282_) );
OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_3278_), .B(_3279_), .C(_3164_), .Y(_3284_) );
NAND3X1 NAND3X1_775 ( .gnd(gnd), .vdd(vdd), .A(_3163_), .B(_3275_), .C(_3276_), .Y(_3285_) );
AOI21X1 AOI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_3284_), .B(_3285_), .C(_3282_), .Y(_3286_) );
OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_3281_), .B(_3286_), .C(_3160_), .Y(_3287_) );
NAND3X1 NAND3X1_776 ( .gnd(gnd), .vdd(vdd), .A(_3282_), .B(_3284_), .C(_3285_), .Y(_3288_) );
NAND3X1 NAND3X1_777 ( .gnd(gnd), .vdd(vdd), .A(_3161_), .B(_3280_), .C(_3277_), .Y(_3289_) );
NAND3X1 NAND3X1_778 ( .gnd(gnd), .vdd(vdd), .A(_2964_), .B(_3288_), .C(_3289_), .Y(_3290_) );
NAND2X1 NAND2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_3290_), .B(_3287_), .Y(_3291_) );
AOI21X1 AOI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_3159_), .B(_3291_), .C(_1639_), .Y(_3292_) );
OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_3159_), .B(_3291_), .C(_3292_), .Y(_3293_) );
XOR2X1 XOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1895_), .B(module_0_W_143_), .Y(_3295_) );
XOR2X1 XOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_3293_), .B(_3295_), .Y(_3296_) );
XOR2X1 XOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_3296_), .B(_2979_), .Y(_3297_) );
NAND2X1 NAND2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_3157_), .B(_3297_), .Y(_3298_) );
INVX1 INVX1_362 ( .gnd(gnd), .vdd(vdd), .A(_3157_), .Y(_3299_) );
XNOR2X1 XNOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_3296_), .B(_2979_), .Y(_3300_) );
AOI21X1 AOI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_3299_), .B(_3300_), .C(_1893_), .Y(_3301_) );
XNOR2X1 XNOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_3783_), .B(module_0_W_159_), .Y(_3302_) );
NAND3X1 NAND3X1_779 ( .gnd(gnd), .vdd(vdd), .A(_3298_), .B(_3302_), .C(_3301_), .Y(_3303_) );
NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_3299_), .B(_3300_), .Y(_3304_) );
OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_3297_), .B(_3157_), .C(_1648_), .Y(_3306_) );
INVX1 INVX1_363 ( .gnd(gnd), .vdd(vdd), .A(_3302_), .Y(_3307_) );
OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .B(_3304_), .C(_3307_), .Y(_3308_) );
NAND2X1 NAND2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_3303_), .B(_3308_), .Y(_3309_) );
XOR2X1 XOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_3309_), .B(_3002_), .Y(_3310_) );
NAND2X1 NAND2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_3156_), .B(_3310_), .Y(_3311_) );
INVX1 INVX1_364 ( .gnd(gnd), .vdd(vdd), .A(_3156_), .Y(_3312_) );
XNOR2X1 XNOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_3309_), .B(_3002_), .Y(_3313_) );
AOI21X1 AOI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_3313_), .C(_1661_), .Y(_3314_) );
XOR2X1 XOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_3794_), .B(module_0_W_175_), .Y(_3315_) );
NAND3X1 NAND3X1_780 ( .gnd(gnd), .vdd(vdd), .A(_3311_), .B(_3315_), .C(_3314_), .Y(_3317_) );
NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_3313_), .Y(_3318_) );
OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_3310_), .B(_3156_), .C(_1722_), .Y(_3319_) );
INVX1 INVX1_365 ( .gnd(gnd), .vdd(vdd), .A(_3315_), .Y(_3320_) );
OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_3319_), .B(_3318_), .C(_3320_), .Y(_3321_) );
NAND2X1 NAND2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_3317_), .B(_3321_), .Y(_3322_) );
XNOR2X1 XNOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_3322_), .B(_3022_), .Y(_3323_) );
NAND2X1 NAND2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_3155_), .B(_3323_), .Y(_3324_) );
XOR2X1 XOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_3322_), .B(_3022_), .Y(_3325_) );
AOI21X1 AOI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_3154_), .B(_3325_), .C(_1671_), .Y(_3326_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(module_0_W_191_), .Y(_3328_) );
NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_191_), .B(_376_), .Y(_3329_) );
NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_3329_), .B(_3328_), .Y(_3330_) );
NAND3X1 NAND3X1_781 ( .gnd(gnd), .vdd(vdd), .A(_3324_), .B(_3330_), .C(_3326_), .Y(_3331_) );
NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_3154_), .B(_3325_), .Y(_3332_) );
OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_3323_), .B(_3155_), .C(_1718_), .Y(_3333_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3328_), .B(_3329_), .C(_3333_), .D(_3332_), .Y(_3334_) );
NAND2X1 NAND2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_3331_), .B(_3334_), .Y(_3335_) );
XOR2X1 XOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_3335_), .B(_3043_), .Y(_3336_) );
NAND2X1 NAND2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_3153_), .B(_3336_), .Y(_3337_) );
INVX1 INVX1_366 ( .gnd(gnd), .vdd(vdd), .A(_3153_), .Y(_3339_) );
XNOR2X1 XNOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_3335_), .B(_3043_), .Y(_3340_) );
AOI21X1 AOI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_3339_), .B(_3340_), .C(_1957_), .Y(_3341_) );
OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_3815_), .B(_3818_), .C(module_0_W_207_), .Y(_3342_) );
INVX1 INVX1_367 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_207_), .Y(_3343_) );
NAND3X1 NAND3X1_782 ( .gnd(gnd), .vdd(vdd), .A(_3343_), .B(_3817_), .C(_3822_), .Y(_3344_) );
NAND2X1 NAND2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_3344_), .B(_3342_), .Y(_3345_) );
INVX1 INVX1_368 ( .gnd(gnd), .vdd(vdd), .A(_3345_), .Y(_3346_) );
NAND3X1 NAND3X1_783 ( .gnd(gnd), .vdd(vdd), .A(_3337_), .B(_3346_), .C(_3341_), .Y(_3347_) );
NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_3339_), .B(_3340_), .Y(_3348_) );
OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(_3153_), .C(_1680_), .Y(_3350_) );
OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_3350_), .B(_3348_), .C(_3345_), .Y(_3351_) );
NAND2X1 NAND2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_3347_), .B(_3351_), .Y(_3352_) );
XOR2X1 XOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_3352_), .B(_3063_), .Y(_3353_) );
XNOR2X1 XNOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_3353_), .B(_3152_), .Y(_3354_) );
OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_3830_), .B(_3833_), .C(module_0_W_223_), .Y(_3355_) );
INVX1 INVX1_369 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_223_), .Y(_3356_) );
NAND2X1 NAND2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_3356_), .B(_3835_), .Y(_3357_) );
NAND2X1 NAND2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_3355_), .B(_3357_), .Y(_3358_) );
NOR3X1 NOR3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_3358_), .B(_1691_), .C(_3354_), .Y(_3359_) );
XOR2X1 XOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_3353_), .B(_3152_), .Y(_3361_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_3357_), .B(_3355_), .Y(_3362_) );
AOI21X1 AOI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_1970_), .B(_3361_), .C(_3362_), .Y(_3363_) );
OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_3359_), .B(_3363_), .C(_3087_), .Y(_3364_) );
INVX1 INVX1_370 ( .gnd(gnd), .vdd(vdd), .A(_3087_), .Y(_3365_) );
NAND3X1 NAND3X1_784 ( .gnd(gnd), .vdd(vdd), .A(_1970_), .B(_3361_), .C(_3362_), .Y(_3366_) );
OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_3354_), .B(_1691_), .C(_3358_), .Y(_3367_) );
NAND3X1 NAND3X1_785 ( .gnd(gnd), .vdd(vdd), .A(_3365_), .B(_3366_), .C(_3367_), .Y(_3368_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_3364_), .B(_3368_), .Y(_3369_) );
NAND2X1 NAND2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_3150_), .B(_3369_), .Y(_3370_) );
INVX1 INVX1_371 ( .gnd(gnd), .vdd(vdd), .A(_3150_), .Y(_3372_) );
NAND2X1 NAND2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_3368_), .B(_3364_), .Y(_3373_) );
AOI21X1 AOI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_3373_), .B(_3372_), .C(_1701_), .Y(_3374_) );
OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_3846_), .B(_3841_), .C(module_0_W_239_), .Y(_3375_) );
INVX1 INVX1_372 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_239_), .Y(_3376_) );
NAND3X1 NAND3X1_786 ( .gnd(gnd), .vdd(vdd), .A(_3376_), .B(_3840_), .C(_3845_), .Y(_3377_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_3375_), .B(_3377_), .Y(_3378_) );
NAND3X1 NAND3X1_787 ( .gnd(gnd), .vdd(vdd), .A(_3370_), .B(_3374_), .C(_3378_), .Y(_3379_) );
NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_3373_), .B(_3372_), .Y(_3380_) );
OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_3150_), .C(_1714_), .Y(_3381_) );
NAND2X1 NAND2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_3377_), .B(_3375_), .Y(_3383_) );
OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_3381_), .B(_3380_), .C(_3383_), .Y(_3384_) );
NAND2X1 NAND2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_3384_), .B(_3379_), .Y(_3385_) );
XNOR2X1 XNOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_3109_), .Y(_3386_) );
NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_3149_), .B(_3386_), .Y(_3387_) );
XOR2X1 XOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_3109_), .Y(_3388_) );
OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_3148_), .C(_1713_), .Y(_3389_) );
OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_3389_), .B(_3387_), .C(_3147_), .Y(_3390_) );
OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_3128_), .B(_3122_), .C(_3388_), .Y(_3391_) );
AOI21X1 AOI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_3149_), .B(_3386_), .C(_1712_), .Y(_3392_) );
NAND3X1 NAND3X1_788 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_255_), .B(_3391_), .C(_3392_), .Y(_3394_) );
NAND3X1 NAND3X1_789 ( .gnd(gnd), .vdd(vdd), .A(_3146_), .B(_3394_), .C(_3390_), .Y(_3395_) );
NAND3X1 NAND3X1_790 ( .gnd(gnd), .vdd(vdd), .A(_3147_), .B(_3391_), .C(_3392_), .Y(_3396_) );
OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_3389_), .B(_3387_), .C(module_0_W_255_), .Y(_3397_) );
NAND3X1 NAND3X1_791 ( .gnd(gnd), .vdd(vdd), .A(_3133_), .B(_3396_), .C(_3397_), .Y(_3398_) );
NAND2X1 NAND2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_3398_), .B(_3395_), .Y(_3399_) );
XNOR2X1 XNOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_3145_), .B(_3399_), .Y(module_0_H_23_) );
INVX1 INVX1_373 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_241_), .Y(_1949_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_0_), .B(module_0_W_16_), .Y(_1960_) );
NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_0_), .B(module_0_W_16_), .Y(_1971_) );
OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_1960_), .B(_1971_), .C(bloque_datos[0]), .Y(_1982_) );
INVX1 INVX1_374 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(_1993_) );
NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_1960_), .Y(_2004_) );
NAND2X1 NAND2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_1993_), .B(_2004_), .Y(_2015_) );
NAND2X1 NAND2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_1982_), .B(_2015_), .Y(_2026_) );
NAND2X1 NAND2X1_428 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf3_), .B(_2026_), .Y(_2037_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_2026_), .B(bloque_datos_16_bF_buf2_), .Y(_2048_) );
NAND2X1 NAND2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_2037_), .B(_2048_), .Y(_2057_) );
NAND2X1 NAND2X1_430 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf4_), .B(_2057_), .Y(_2066_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_2057_), .B(bloque_datos_32_bF_buf3_), .Y(_2076_) );
NAND2X1 NAND2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_2066_), .B(_2076_), .Y(_2087_) );
NAND2X1 NAND2X1_432 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_48_bF_buf4_), .B(_2087_), .Y(_2098_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_2087_), .B(bloque_datos_48_bF_buf3_), .Y(_2109_) );
NAND2X1 NAND2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_2098_), .B(_2109_), .Y(_2120_) );
NAND2X1 NAND2X1_434 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_64_bF_buf4_), .B(_2120_), .Y(_2131_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_2120_), .B(bloque_datos_64_bF_buf3_), .Y(_2142_) );
NAND2X1 NAND2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_2131_), .B(_2142_), .Y(_2153_) );
NAND2X1 NAND2X1_436 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf5_), .B(_2153_), .Y(_2164_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_2153_), .B(bloque_datos_80_bF_buf4_), .Y(_2175_) );
NAND2X1 NAND2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_2164_), .B(_2175_), .Y(_2186_) );
NAND2X1 NAND2X1_438 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_128_), .B(_2186_), .Y(_2197_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(module_0_W_128_), .Y(_2208_) );
NAND2X1 NAND2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_2197_), .B(_2208_), .Y(_2219_) );
NAND2X1 NAND2X1_440 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_144_), .B(_2219_), .Y(_2230_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_2219_), .B(module_0_W_144_), .Y(_2241_) );
NAND2X1 NAND2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_2230_), .B(_2241_), .Y(_2252_) );
NAND2X1 NAND2X1_442 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_160_), .B(_2252_), .Y(_2263_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_2252_), .B(module_0_W_160_), .Y(_2274_) );
NAND2X1 NAND2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_2263_), .B(_2274_), .Y(_2285_) );
NAND2X1 NAND2X1_444 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_176_), .B(_2285_), .Y(_2296_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_2285_), .B(module_0_W_176_), .Y(_2307_) );
NAND2X1 NAND2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_2296_), .B(_2307_), .Y(_2318_) );
NAND2X1 NAND2X1_446 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_192_), .B(_2318_), .Y(_2329_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_2318_), .B(module_0_W_192_), .Y(_2340_) );
NAND2X1 NAND2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_2329_), .B(_2340_), .Y(_2351_) );
NAND2X1 NAND2X1_448 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_208_), .B(_2351_), .Y(_2362_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_2351_), .B(module_0_W_208_), .Y(_2373_) );
NAND2X1 NAND2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_2362_), .B(_2373_), .Y(_2384_) );
INVX2 INVX2_72 ( .gnd(gnd), .vdd(vdd), .A(_2384_), .Y(_2395_) );
NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_224_), .B(_2395_), .Y(_2406_) );
INVX1 INVX1_375 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_225_), .Y(_2417_) );
INVX2 INVX2_73 ( .gnd(gnd), .vdd(vdd), .A(_2351_), .Y(_2428_) );
NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_208_), .B(_2428_), .Y(_2439_) );
INVX2 INVX2_74 ( .gnd(gnd), .vdd(vdd), .A(_2318_), .Y(_2449_) );
NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_192_), .B(_2449_), .Y(_2460_) );
INVX1 INVX1_376 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_193_), .Y(_2471_) );
INVX2 INVX2_75 ( .gnd(gnd), .vdd(vdd), .A(_2285_), .Y(_2482_) );
NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_176_), .B(_2482_), .Y(_2493_) );
INVX2 INVX2_76 ( .gnd(gnd), .vdd(vdd), .A(_2252_), .Y(_2504_) );
NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_160_), .B(_2504_), .Y(_2515_) );
INVX1 INVX1_377 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_161_), .Y(_2526_) );
INVX2 INVX2_77 ( .gnd(gnd), .vdd(vdd), .A(_2219_), .Y(_2537_) );
NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_144_), .B(_2537_), .Y(_2548_) );
INVX1 INVX1_378 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_145_), .Y(_2559_) );
INVX2 INVX2_78 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .Y(_2570_) );
NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_128_), .B(_2570_), .Y(_2581_) );
INVX2 INVX2_79 ( .gnd(gnd), .vdd(vdd), .A(_2153_), .Y(_2592_) );
NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf3_), .B(_2592_), .Y(_2603_) );
AOI21X1 AOI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_2098_), .B(_2109_), .C(bloque_datos_64_bF_buf2_), .Y(_2614_) );
AOI21X1 AOI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_2066_), .B(_2076_), .C(bloque_datos_48_bF_buf2_), .Y(_2625_) );
INVX1 INVX1_379 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_49_bF_buf3_), .Y(_2636_) );
AOI21X1 AOI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_2037_), .B(_2048_), .C(bloque_datos_32_bF_buf2_), .Y(_2647_) );
INVX1 INVX1_380 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf3_), .Y(_2658_) );
AOI21X1 AOI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_1982_), .B(_2015_), .C(bloque_datos_16_bF_buf1_), .Y(_2669_) );
OAI21X1 OAI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_1960_), .B(_1971_), .C(_1993_), .Y(_2680_) );
INVX1 INVX1_381 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(_2691_) );
INVX2 INVX2_80 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_0_), .Y(_2702_) );
NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_16_), .B(_2702_), .Y(_2713_) );
NAND2X1 NAND2X1_450 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_0_), .B(module_0_W_1_), .Y(_2724_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_0_), .B(module_0_W_1_), .Y(_2735_) );
AOI21X1 AOI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_2724_), .B(_2735_), .C(module_0_W_17_), .Y(_2746_) );
INVX1 INVX1_382 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_17_), .Y(_2757_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_0_), .B(module_0_W_1_), .Y(_2768_) );
NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_0_), .B(module_0_W_1_), .Y(_2779_) );
NOR3X1 NOR3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_2757_), .B(_2779_), .C(_2768_), .Y(_2790_) );
OAI21X1 OAI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_2790_), .B(_2746_), .C(_2713_), .Y(_2801_) );
INVX1 INVX1_383 ( .gnd(gnd), .vdd(vdd), .A(_2713_), .Y(_2811_) );
OAI21X1 OAI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .B(_2779_), .C(_2757_), .Y(_2822_) );
NAND3X1 NAND3X1_792 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_17_), .B(_2724_), .C(_2735_), .Y(_2833_) );
NAND3X1 NAND3X1_793 ( .gnd(gnd), .vdd(vdd), .A(_2822_), .B(_2833_), .C(_2811_), .Y(_2844_) );
NAND2X1 NAND2X1_451 ( .gnd(gnd), .vdd(vdd), .A(_2844_), .B(_2801_), .Y(_2855_) );
NAND2X1 NAND2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_2691_), .B(_2855_), .Y(_2866_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_2855_), .B(_2691_), .Y(_2877_) );
NAND2X1 NAND2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_2866_), .B(_2877_), .Y(_2888_) );
XNOR2X1 XNOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_2888_), .B(_2680_), .Y(_2899_) );
XNOR2X1 XNOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_2899_), .B(bloque_datos[17]), .Y(_2910_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_2910_), .B(_2669_), .Y(_2921_) );
NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_2669_), .B(_2910_), .Y(_2932_) );
OAI21X1 OAI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_2921_), .B(_2932_), .C(_2658_), .Y(_2943_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_2921_), .B(_2932_), .Y(_2954_) );
NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .B(_2954_), .Y(_2965_) );
INVX1 INVX1_384 ( .gnd(gnd), .vdd(vdd), .A(_2965_), .Y(_2976_) );
NAND2X1 NAND2X1_454 ( .gnd(gnd), .vdd(vdd), .A(_2943_), .B(_2976_), .Y(_2987_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_2987_), .B(_2647_), .Y(_2998_) );
NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_2647_), .B(_2987_), .Y(_3009_) );
OAI21X1 OAI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_2998_), .B(_3009_), .C(_2636_), .Y(_3020_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_2998_), .B(_3009_), .Y(_3031_) );
NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_2636_), .B(_3031_), .Y(_3042_) );
INVX1 INVX1_385 ( .gnd(gnd), .vdd(vdd), .A(_3042_), .Y(_3053_) );
NAND2X1 NAND2X1_455 ( .gnd(gnd), .vdd(vdd), .A(_3020_), .B(_3053_), .Y(_3064_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_3064_), .B(_2625_), .Y(_3075_) );
NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .B(_3064_), .Y(_3086_) );
NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_3086_), .B(_3075_), .Y(_3097_) );
XNOR2X1 XNOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_3097_), .B(bloque_datos_65_bF_buf3_), .Y(_3108_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_3108_), .B(_2614_), .Y(_3119_) );
NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_2614_), .B(_3108_), .Y(_3130_) );
NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_3130_), .B(_3119_), .Y(_3141_) );
NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf4_), .B(_3141_), .Y(_3151_) );
INVX1 INVX1_386 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf3_), .Y(_3162_) );
INVX1 INVX1_387 ( .gnd(gnd), .vdd(vdd), .A(_3141_), .Y(_3173_) );
NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_3162_), .B(_3173_), .Y(_3184_) );
OAI21X1 OAI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_3184_), .B(_3151_), .C(_2603_), .Y(_3195_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_3184_), .B(_3151_), .Y(_3206_) );
NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_2603_), .B(_3206_), .Y(_3217_) );
INVX2 INVX2_81 ( .gnd(gnd), .vdd(vdd), .A(_3217_), .Y(_3228_) );
NAND2X1 NAND2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_3195_), .B(_3228_), .Y(_3239_) );
INVX2 INVX2_82 ( .gnd(gnd), .vdd(vdd), .A(_3239_), .Y(_3250_) );
NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_129_), .B(_3250_), .Y(_3261_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_3250_), .B(module_0_W_129_), .Y(_3272_) );
OAI21X1 OAI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_3272_), .B(_3261_), .C(_2581_), .Y(_3283_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_3272_), .B(_3261_), .Y(_3294_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_3294_), .B(_2581_), .Y(_3305_) );
NAND2X1 NAND2X1_457 ( .gnd(gnd), .vdd(vdd), .A(_3283_), .B(_3305_), .Y(_3316_) );
NAND2X1 NAND2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2559_), .B(_3316_), .Y(_3327_) );
NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_2559_), .B(_3316_), .Y(_3338_) );
INVX1 INVX1_388 ( .gnd(gnd), .vdd(vdd), .A(_3338_), .Y(_3349_) );
NAND2X1 NAND2X1_459 ( .gnd(gnd), .vdd(vdd), .A(_3327_), .B(_3349_), .Y(_3360_) );
NAND2X1 NAND2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_2548_), .B(_3360_), .Y(_3371_) );
NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_2548_), .B(_3360_), .Y(_3382_) );
INVX1 INVX1_389 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .Y(_3393_) );
NAND2X1 NAND2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_3371_), .B(_3393_), .Y(_3400_) );
NAND2X1 NAND2X1_462 ( .gnd(gnd), .vdd(vdd), .A(_2526_), .B(_3400_), .Y(_3401_) );
NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_2526_), .B(_3400_), .Y(_3402_) );
INVX1 INVX1_390 ( .gnd(gnd), .vdd(vdd), .A(_3402_), .Y(_3403_) );
NAND2X1 NAND2X1_463 ( .gnd(gnd), .vdd(vdd), .A(_3401_), .B(_3403_), .Y(_3404_) );
NAND2X1 NAND2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_2515_), .B(_3404_), .Y(_3405_) );
NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_2515_), .B(_3404_), .Y(_3406_) );
INVX1 INVX1_391 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .Y(_3407_) );
NAND2X1 NAND2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_3405_), .B(_3407_), .Y(_3408_) );
INVX2 INVX2_83 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .Y(_3409_) );
NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_177_), .B(_3409_), .Y(_3410_) );
NAND2X1 NAND2X1_466 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_177_), .B(_3409_), .Y(_3411_) );
INVX2 INVX2_84 ( .gnd(gnd), .vdd(vdd), .A(_3411_), .Y(_3412_) );
OAI21X1 OAI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_3412_), .B(_3410_), .C(_2493_), .Y(_3413_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_3412_), .B(_3410_), .Y(_3414_) );
NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_2493_), .B(_3414_), .Y(_3415_) );
INVX1 INVX1_392 ( .gnd(gnd), .vdd(vdd), .A(_3415_), .Y(_3416_) );
NAND2X1 NAND2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_3413_), .B(_3416_), .Y(_3417_) );
NAND2X1 NAND2X1_468 ( .gnd(gnd), .vdd(vdd), .A(_2471_), .B(_3417_), .Y(_3418_) );
NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_2471_), .B(_3417_), .Y(_3419_) );
INVX1 INVX1_393 ( .gnd(gnd), .vdd(vdd), .A(_3419_), .Y(_3420_) );
NAND2X1 NAND2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_3418_), .B(_3420_), .Y(_3421_) );
NAND2X1 NAND2X1_470 ( .gnd(gnd), .vdd(vdd), .A(_2460_), .B(_3421_), .Y(_3422_) );
NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_2460_), .B(_3421_), .Y(_3423_) );
INVX1 INVX1_394 ( .gnd(gnd), .vdd(vdd), .A(_3423_), .Y(_3424_) );
NAND2X1 NAND2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_3422_), .B(_3424_), .Y(_3425_) );
INVX2 INVX2_85 ( .gnd(gnd), .vdd(vdd), .A(_3425_), .Y(_3426_) );
NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_209_), .B(_3426_), .Y(_3427_) );
NAND2X1 NAND2X1_472 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_209_), .B(_3426_), .Y(_3428_) );
INVX2 INVX2_86 ( .gnd(gnd), .vdd(vdd), .A(_3428_), .Y(_3429_) );
OAI21X1 OAI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_3429_), .B(_3427_), .C(_2439_), .Y(_3430_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_3429_), .B(_3427_), .Y(_3431_) );
NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_2439_), .B(_3431_), .Y(_3432_) );
INVX2 INVX2_87 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3433_) );
NAND2X1 NAND2X1_473 ( .gnd(gnd), .vdd(vdd), .A(_3430_), .B(_3433_), .Y(_3434_) );
NAND2X1 NAND2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_2417_), .B(_3434_), .Y(_3435_) );
NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_2417_), .B(_3434_), .Y(_3436_) );
INVX1 INVX1_395 ( .gnd(gnd), .vdd(vdd), .A(_3436_), .Y(_3437_) );
NAND2X1 NAND2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_3435_), .B(_3437_), .Y(_3438_) );
NAND2X1 NAND2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_2406_), .B(_3438_), .Y(_3439_) );
NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_2406_), .B(_3438_), .Y(_3440_) );
INVX1 INVX1_396 ( .gnd(gnd), .vdd(vdd), .A(_3440_), .Y(_3441_) );
NAND2X1 NAND2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_3439_), .B(_3441_), .Y(_3442_) );
NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1949_), .B(_3442_), .Y(_3443_) );
INVX1 INVX1_397 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_242_), .Y(_3444_) );
INVX1 INVX1_398 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_194_), .Y(_3445_) );
INVX1 INVX1_399 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_178_), .Y(_3446_) );
INVX1 INVX1_400 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_162_), .Y(_3447_) );
NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_2581_), .B(_3294_), .Y(_3448_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_3097_), .B(bloque_datos_65_bF_buf2_), .Y(_3449_) );
INVX1 INVX1_401 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf4_), .Y(_3450_) );
INVX1 INVX1_402 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf4_), .Y(_3451_) );
INVX1 INVX1_403 ( .gnd(gnd), .vdd(vdd), .A(_2932_), .Y(_3452_) );
NAND2X1 NAND2X1_478 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .B(_2899_), .Y(_3453_) );
INVX1 INVX1_404 ( .gnd(gnd), .vdd(vdd), .A(_2680_), .Y(_3454_) );
NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_3454_), .B(_2888_), .Y(_3455_) );
INVX1 INVX1_405 ( .gnd(gnd), .vdd(vdd), .A(_2877_), .Y(_3456_) );
INVX1 INVX1_406 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf3_), .Y(_3457_) );
INVX1 INVX1_407 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_18_), .Y(_3458_) );
NAND3X1 NAND3X1_794 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_2_), .B(module_0_W_0_), .C(module_0_W_1_), .Y(_3459_) );
INVX2 INVX2_88 ( .gnd(gnd), .vdd(vdd), .A(_3459_), .Y(_3460_) );
AOI21X1 AOI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_0_), .B(module_0_W_1_), .C(module_0_W_2_), .Y(_3461_) );
OAI21X1 OAI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_3460_), .B(_3461_), .C(_3458_), .Y(_3462_) );
INVX2 INVX2_89 ( .gnd(gnd), .vdd(vdd), .A(_3461_), .Y(_3463_) );
NAND3X1 NAND3X1_795 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_18_), .B(_3459_), .C(_3463_), .Y(_3464_) );
NAND3X1 NAND3X1_796 ( .gnd(gnd), .vdd(vdd), .A(_2790_), .B(_3464_), .C(_3462_), .Y(_3465_) );
AOI21X1 AOI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_3459_), .B(_3463_), .C(module_0_W_18_), .Y(_3466_) );
NOR3X1 NOR3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_3458_), .B(_3461_), .C(_3460_), .Y(_3467_) );
OAI21X1 OAI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_3467_), .B(_3466_), .C(_2833_), .Y(_3468_) );
NAND2X1 NAND2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_3465_), .B(_3468_), .Y(_3469_) );
NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_2844_), .B(_3469_), .Y(_3470_) );
INVX1 INVX1_408 ( .gnd(gnd), .vdd(vdd), .A(_2844_), .Y(_3471_) );
AOI21X1 AOI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_3465_), .B(_3468_), .C(_3471_), .Y(_3472_) );
OAI21X1 OAI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_3470_), .B(_3472_), .C(_3457_), .Y(_3473_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_3469_), .B(_2844_), .Y(_3474_) );
INVX1 INVX1_409 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .Y(_3475_) );
NAND3X1 NAND3X1_797 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf2_), .B(_3475_), .C(_3474_), .Y(_3476_) );
NAND3X1 NAND3X1_798 ( .gnd(gnd), .vdd(vdd), .A(_3456_), .B(_3473_), .C(_3476_), .Y(_3477_) );
AOI21X1 AOI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_3475_), .B(_3474_), .C(bloque_datos_2_bF_buf1_), .Y(_3478_) );
NOR3X1 NOR3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_3457_), .B(_3472_), .C(_3470_), .Y(_3479_) );
OAI21X1 OAI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_3478_), .B(_3479_), .C(_2877_), .Y(_3480_) );
NAND3X1 NAND3X1_799 ( .gnd(gnd), .vdd(vdd), .A(_3455_), .B(_3477_), .C(_3480_), .Y(_3481_) );
AOI21X1 AOI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_3477_), .B(_3480_), .C(_3455_), .Y(_3482_) );
INVX1 INVX1_410 ( .gnd(gnd), .vdd(vdd), .A(_3482_), .Y(_3483_) );
AOI21X1 AOI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_3481_), .B(_3483_), .C(bloque_datos[18]), .Y(_3484_) );
INVX1 INVX1_411 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .Y(_3485_) );
INVX1 INVX1_412 ( .gnd(gnd), .vdd(vdd), .A(_3455_), .Y(_3486_) );
NOR3X1 NOR3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_3479_), .B(_2877_), .C(_3478_), .Y(_3487_) );
AOI21X1 AOI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .B(_3476_), .C(_3456_), .Y(_3488_) );
NOR3X1 NOR3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_3486_), .B(_3488_), .C(_3487_), .Y(_3489_) );
NOR3X1 NOR3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_3485_), .B(_3482_), .C(_3489_), .Y(_3490_) );
NOR3X1 NOR3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_3453_), .B(_3490_), .C(_3484_), .Y(_3491_) );
INVX1 INVX1_413 ( .gnd(gnd), .vdd(vdd), .A(_3453_), .Y(_3492_) );
OAI21X1 OAI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_3489_), .B(_3482_), .C(_3485_), .Y(_3493_) );
INVX2 INVX2_90 ( .gnd(gnd), .vdd(vdd), .A(_3490_), .Y(_3494_) );
AOI21X1 AOI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_3493_), .B(_3494_), .C(_3492_), .Y(_3495_) );
NOR3X1 NOR3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_3452_), .B(_3491_), .C(_3495_), .Y(_3496_) );
NAND3X1 NAND3X1_800 ( .gnd(gnd), .vdd(vdd), .A(_3492_), .B(_3493_), .C(_3494_), .Y(_3497_) );
OAI21X1 OAI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_3484_), .B(_3490_), .C(_3453_), .Y(_3498_) );
AOI21X1 AOI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_3497_), .C(_2932_), .Y(_3499_) );
OAI21X1 OAI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_3496_), .B(_3499_), .C(_3451_), .Y(_3500_) );
NAND3X1 NAND3X1_801 ( .gnd(gnd), .vdd(vdd), .A(_2932_), .B(_3498_), .C(_3497_), .Y(_3501_) );
OAI21X1 OAI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_3495_), .B(_3491_), .C(_3452_), .Y(_3502_) );
NAND3X1 NAND3X1_802 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf3_), .B(_3501_), .C(_3502_), .Y(_3503_) );
NAND3X1 NAND3X1_803 ( .gnd(gnd), .vdd(vdd), .A(_2965_), .B(_3503_), .C(_3500_), .Y(_3504_) );
AOI21X1 AOI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_3501_), .B(_3502_), .C(bloque_datos_34_bF_buf2_), .Y(_3505_) );
NOR3X1 NOR3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .B(_3499_), .C(_3496_), .Y(_3506_) );
OAI21X1 OAI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_3506_), .B(_3505_), .C(_2976_), .Y(_3507_) );
NAND3X1 NAND3X1_804 ( .gnd(gnd), .vdd(vdd), .A(_3009_), .B(_3504_), .C(_3507_), .Y(_3508_) );
AOI21X1 AOI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_3504_), .B(_3507_), .C(_3009_), .Y(_3509_) );
INVX1 INVX1_414 ( .gnd(gnd), .vdd(vdd), .A(_3509_), .Y(_3510_) );
AOI21X1 AOI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_3510_), .C(bloque_datos_50_bF_buf3_), .Y(_3511_) );
INVX1 INVX1_415 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_50_bF_buf2_), .Y(_3512_) );
INVX1 INVX1_416 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .Y(_3513_) );
NOR3X1 NOR3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_3512_), .B(_3509_), .C(_3513_), .Y(_3514_) );
NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_3511_), .B(_3514_), .Y(_3515_) );
NAND2X1 NAND2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_3042_), .B(_3515_), .Y(_3516_) );
OAI21X1 OAI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_3514_), .B(_3511_), .C(_3053_), .Y(_3517_) );
NAND3X1 NAND3X1_805 ( .gnd(gnd), .vdd(vdd), .A(_3086_), .B(_3517_), .C(_3516_), .Y(_3518_) );
INVX2 INVX2_91 ( .gnd(gnd), .vdd(vdd), .A(_3518_), .Y(_3519_) );
AOI21X1 AOI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_3517_), .B(_3516_), .C(_3086_), .Y(_3520_) );
OAI21X1 OAI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_3519_), .B(_3520_), .C(_3450_), .Y(_3521_) );
INVX1 INVX1_417 ( .gnd(gnd), .vdd(vdd), .A(_3086_), .Y(_3522_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_3515_), .B(_3042_), .Y(_3523_) );
INVX1 INVX1_418 ( .gnd(gnd), .vdd(vdd), .A(_3517_), .Y(_3524_) );
OAI21X1 OAI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_3523_), .B(_3524_), .C(_3522_), .Y(_3525_) );
NAND3X1 NAND3X1_806 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf3_), .B(_3518_), .C(_3525_), .Y(_3526_) );
NAND3X1 NAND3X1_807 ( .gnd(gnd), .vdd(vdd), .A(_3449_), .B(_3526_), .C(_3521_), .Y(_3527_) );
INVX1 INVX1_419 ( .gnd(gnd), .vdd(vdd), .A(_3449_), .Y(_3528_) );
AOI21X1 AOI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_3518_), .B(_3525_), .C(bloque_datos_66_bF_buf2_), .Y(_3529_) );
NOR3X1 NOR3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_3450_), .B(_3520_), .C(_3519_), .Y(_3530_) );
OAI21X1 OAI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(_3529_), .C(_3528_), .Y(_3531_) );
NAND3X1 NAND3X1_808 ( .gnd(gnd), .vdd(vdd), .A(_3130_), .B(_3527_), .C(_3531_), .Y(_3532_) );
INVX2 INVX2_92 ( .gnd(gnd), .vdd(vdd), .A(_3130_), .Y(_3533_) );
NOR3X1 NOR3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_3528_), .B(_3529_), .C(_3530_), .Y(_3534_) );
AOI21X1 AOI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_3526_), .B(_3521_), .C(_3449_), .Y(_3535_) );
OAI21X1 OAI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_3534_), .B(_3535_), .C(_3533_), .Y(_3536_) );
AOI21X1 AOI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_3536_), .C(bloque_datos_82_bF_buf4_), .Y(_3537_) );
INVX1 INVX1_420 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf3_), .Y(_3538_) );
NOR3X1 NOR3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_3533_), .B(_3535_), .C(_3534_), .Y(_3539_) );
AOI21X1 AOI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_3527_), .B(_3531_), .C(_3130_), .Y(_3540_) );
NOR3X1 NOR3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_3538_), .B(_3540_), .C(_3539_), .Y(_3541_) );
NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_3537_), .B(_3541_), .Y(_3542_) );
NAND2X1 NAND2X1_481 ( .gnd(gnd), .vdd(vdd), .A(_3184_), .B(_3542_), .Y(_3543_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_3162_), .B(_3173_), .C(_3541_), .D(_3537_), .Y(_3544_) );
NAND3X1 NAND3X1_809 ( .gnd(gnd), .vdd(vdd), .A(_3217_), .B(_3544_), .C(_3543_), .Y(_3545_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_3542_), .B(_3184_), .Y(_3546_) );
INVX2 INVX2_93 ( .gnd(gnd), .vdd(vdd), .A(_3544_), .Y(_3547_) );
OAI21X1 OAI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_3546_), .B(_3547_), .C(_3228_), .Y(_3548_) );
AOI21X1 AOI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_3545_), .B(_3548_), .C(module_0_W_130_), .Y(_3549_) );
INVX1 INVX1_421 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_130_), .Y(_3550_) );
NOR3X1 NOR3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_3547_), .B(_3228_), .C(_3546_), .Y(_3551_) );
AOI21X1 AOI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_3544_), .B(_3543_), .C(_3217_), .Y(_3552_) );
NOR3X1 NOR3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_3550_), .B(_3552_), .C(_3551_), .Y(_3553_) );
NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_3549_), .B(_3553_), .Y(_3554_) );
NAND2X1 NAND2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_3272_), .B(_3554_), .Y(_3555_) );
NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_3272_), .B(_3554_), .Y(_3556_) );
INVX1 INVX1_422 ( .gnd(gnd), .vdd(vdd), .A(_3556_), .Y(_3557_) );
NAND3X1 NAND3X1_810 ( .gnd(gnd), .vdd(vdd), .A(_3448_), .B(_3555_), .C(_3557_), .Y(_3558_) );
INVX1 INVX1_423 ( .gnd(gnd), .vdd(vdd), .A(_3555_), .Y(_3559_) );
OAI21X1 OAI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_3559_), .B(_3556_), .C(_3305_), .Y(_3560_) );
AOI21X1 AOI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_3560_), .B(_3558_), .C(module_0_W_146_), .Y(_3561_) );
INVX1 INVX1_424 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_146_), .Y(_3562_) );
NOR3X1 NOR3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_3305_), .B(_3556_), .C(_3559_), .Y(_3563_) );
AOI21X1 AOI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_3555_), .B(_3557_), .C(_3448_), .Y(_3564_) );
NOR3X1 NOR3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_3563_), .B(_3562_), .C(_3564_), .Y(_3565_) );
NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_3561_), .B(_3565_), .Y(_3566_) );
NAND2X1 NAND2X1_483 ( .gnd(gnd), .vdd(vdd), .A(_3338_), .B(_3566_), .Y(_3567_) );
OAI21X1 OAI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_3565_), .B(_3561_), .C(_3349_), .Y(_3568_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_3567_), .B(_3568_), .Y(_3569_) );
NAND2X1 NAND2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .B(_3569_), .Y(_3570_) );
INVX1 INVX1_425 ( .gnd(gnd), .vdd(vdd), .A(_3570_), .Y(_3571_) );
NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .B(_3569_), .Y(_3572_) );
OAI21X1 OAI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_3571_), .B(_3572_), .C(_3447_), .Y(_3573_) );
NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_3572_), .B(_3571_), .Y(_3574_) );
NAND2X1 NAND2X1_485 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_162_), .B(_3574_), .Y(_3575_) );
NAND3X1 NAND3X1_811 ( .gnd(gnd), .vdd(vdd), .A(_3402_), .B(_3573_), .C(_3575_), .Y(_3576_) );
INVX1 INVX1_426 ( .gnd(gnd), .vdd(vdd), .A(_3573_), .Y(_3577_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .B(module_0_W_162_), .Y(_3578_) );
OAI21X1 OAI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(_3577_), .C(_3403_), .Y(_3579_) );
NAND3X1 NAND3X1_812 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .B(_3576_), .C(_3579_), .Y(_3580_) );
INVX2 INVX2_94 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .Y(_3581_) );
AOI21X1 AOI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_3576_), .B(_3579_), .C(_3406_), .Y(_3582_) );
OAI21X1 OAI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_3581_), .B(_3582_), .C(_3446_), .Y(_3583_) );
NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_3582_), .B(_3581_), .Y(_3584_) );
NAND2X1 NAND2X1_486 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_178_), .B(_3584_), .Y(_3585_) );
NAND3X1 NAND3X1_813 ( .gnd(gnd), .vdd(vdd), .A(_3412_), .B(_3583_), .C(_3585_), .Y(_3586_) );
INVX1 INVX1_427 ( .gnd(gnd), .vdd(vdd), .A(_3583_), .Y(_3587_) );
INVX1 INVX1_428 ( .gnd(gnd), .vdd(vdd), .A(_3585_), .Y(_3588_) );
OAI21X1 OAI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_3588_), .B(_3587_), .C(_3411_), .Y(_3589_) );
NAND3X1 NAND3X1_814 ( .gnd(gnd), .vdd(vdd), .A(_3415_), .B(_3586_), .C(_3589_), .Y(_3590_) );
INVX2 INVX2_95 ( .gnd(gnd), .vdd(vdd), .A(_3590_), .Y(_3591_) );
AOI21X1 AOI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_3586_), .B(_3589_), .C(_3415_), .Y(_3592_) );
OAI21X1 OAI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_3591_), .B(_3592_), .C(_3445_), .Y(_3593_) );
INVX1 INVX1_429 ( .gnd(gnd), .vdd(vdd), .A(_3593_), .Y(_3594_) );
NOR3X1 NOR3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_3445_), .B(_3592_), .C(_3591_), .Y(_3595_) );
NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_3595_), .B(_3594_), .Y(_3596_) );
NAND2X1 NAND2X1_487 ( .gnd(gnd), .vdd(vdd), .A(_3419_), .B(_3596_), .Y(_3597_) );
OAI21X1 OAI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_3594_), .B(_3595_), .C(_3420_), .Y(_3598_) );
NAND3X1 NAND3X1_815 ( .gnd(gnd), .vdd(vdd), .A(_3423_), .B(_3598_), .C(_3597_), .Y(_3599_) );
INVX2 INVX2_96 ( .gnd(gnd), .vdd(vdd), .A(_3599_), .Y(_3600_) );
AOI21X1 AOI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_3598_), .B(_3597_), .C(_3423_), .Y(_3601_) );
NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_3601_), .B(_3600_), .Y(_3602_) );
NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_210_), .B(_3602_), .Y(_3603_) );
INVX1 INVX1_430 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_210_), .Y(_3604_) );
NOR3X1 NOR3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_3604_), .B(_3601_), .C(_3600_), .Y(_3605_) );
NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_3605_), .B(_3603_), .Y(_3606_) );
NAND2X1 NAND2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_3429_), .B(_3606_), .Y(_3607_) );
INVX1 INVX1_431 ( .gnd(gnd), .vdd(vdd), .A(_3607_), .Y(_3608_) );
OAI21X1 OAI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_3603_), .B(_3605_), .C(_3428_), .Y(_3609_) );
INVX2 INVX2_97 ( .gnd(gnd), .vdd(vdd), .A(_3609_), .Y(_3610_) );
NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_3610_), .B(_3608_), .Y(_3611_) );
NAND2X1 NAND2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .B(_3611_), .Y(_3612_) );
OAI21X1 OAI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_3608_), .B(_3610_), .C(_3433_), .Y(_3613_) );
AOI21X1 AOI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_3613_), .B(_3612_), .C(module_0_W_226_), .Y(_3614_) );
INVX1 INVX1_432 ( .gnd(gnd), .vdd(vdd), .A(_3614_), .Y(_3615_) );
NAND3X1 NAND3X1_816 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_226_), .B(_3613_), .C(_3612_), .Y(_3616_) );
NAND3X1 NAND3X1_817 ( .gnd(gnd), .vdd(vdd), .A(_3436_), .B(_3616_), .C(_3615_), .Y(_3617_) );
INVX2 INVX2_98 ( .gnd(gnd), .vdd(vdd), .A(_3616_), .Y(_3618_) );
OAI21X1 OAI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_3618_), .B(_3614_), .C(_3437_), .Y(_3619_) );
NAND3X1 NAND3X1_818 ( .gnd(gnd), .vdd(vdd), .A(_3440_), .B(_3619_), .C(_3617_), .Y(_3620_) );
INVX1 INVX1_433 ( .gnd(gnd), .vdd(vdd), .A(_3620_), .Y(_3621_) );
AOI21X1 AOI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_3619_), .B(_3617_), .C(_3440_), .Y(_3622_) );
OAI21X1 OAI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_3621_), .B(_3622_), .C(_3444_), .Y(_3623_) );
NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_3622_), .B(_3621_), .Y(_3624_) );
NAND2X1 NAND2X1_490 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_242_), .B(_3624_), .Y(_3625_) );
NAND3X1 NAND3X1_819 ( .gnd(gnd), .vdd(vdd), .A(_3443_), .B(_3623_), .C(_3625_), .Y(_3626_) );
NAND2X1 NAND2X1_491 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_224_), .B(_2384_), .Y(_3627_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_2384_), .B(module_0_W_224_), .Y(_3628_) );
NAND2X1 NAND2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_3627_), .B(_3628_), .Y(_3629_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(_3629_), .Y(_3630_) );
INVX2 INVX2_99 ( .gnd(gnd), .vdd(vdd), .A(_3442_), .Y(_3631_) );
NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_241_), .B(_3631_), .Y(_3632_) );
NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_3443_), .B(_3632_), .Y(_3633_) );
OAI21X1 OAI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_240_), .B(_3630_), .C(_3633_), .Y(_3634_) );
INVX1 INVX1_434 ( .gnd(gnd), .vdd(vdd), .A(_3443_), .Y(_3635_) );
INVX1 INVX1_435 ( .gnd(gnd), .vdd(vdd), .A(_3623_), .Y(_3636_) );
INVX1 INVX1_436 ( .gnd(gnd), .vdd(vdd), .A(_3625_), .Y(_3637_) );
OAI21X1 OAI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_3637_), .B(_3636_), .C(_3635_), .Y(_3638_) );
INVX1 INVX1_437 ( .gnd(gnd), .vdd(vdd), .A(_3638_), .Y(_3639_) );
OAI21X1 OAI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_3639_), .B(_3634_), .C(_3626_), .Y(_3640_) );
INVX1 INVX1_438 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_243_), .Y(_3641_) );
NAND2X1 NAND2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(_3620_), .Y(_3642_) );
INVX1 INVX1_439 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_227_), .Y(_3643_) );
OAI21X1 OAI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .B(_3610_), .C(_3607_), .Y(_3644_) );
INVX1 INVX1_440 ( .gnd(gnd), .vdd(vdd), .A(_3605_), .Y(_3645_) );
INVX1 INVX1_441 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_211_), .Y(_3646_) );
INVX1 INVX1_442 ( .gnd(gnd), .vdd(vdd), .A(_3597_), .Y(_3647_) );
AOI21X1 AOI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_3423_), .B(_3598_), .C(_3647_), .Y(_3648_) );
INVX1 INVX1_443 ( .gnd(gnd), .vdd(vdd), .A(_3595_), .Y(_3649_) );
INVX1 INVX1_444 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_195_), .Y(_3650_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_3590_), .B(_3586_), .Y(_3651_) );
INVX1 INVX1_445 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_179_), .Y(_3652_) );
INVX1 INVX1_446 ( .gnd(gnd), .vdd(vdd), .A(_3576_), .Y(_3653_) );
INVX1 INVX1_447 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_163_), .Y(_3654_) );
INVX1 INVX1_448 ( .gnd(gnd), .vdd(vdd), .A(_3568_), .Y(_3655_) );
OAI21X1 OAI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .B(_3655_), .C(_3567_), .Y(_3656_) );
INVX1 INVX1_449 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_147_), .Y(_3657_) );
OAI21X1 OAI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_3305_), .B(_3556_), .C(_3555_), .Y(_3658_) );
INVX1 INVX1_450 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_131_), .Y(_3659_) );
OAI21X1 OAI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_3228_), .B(_3547_), .C(_3543_), .Y(_3660_) );
OAI21X1 OAI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_3535_), .B(_3533_), .C(_3527_), .Y(_3661_) );
OAI21X1 OAI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_3524_), .B(_3522_), .C(_3516_), .Y(_3662_) );
INVX1 INVX1_451 ( .gnd(gnd), .vdd(vdd), .A(_3514_), .Y(_3663_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_3504_), .Y(_3664_) );
AOI21X1 AOI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_2932_), .C(_3491_), .Y(_3665_) );
INVX2 INVX2_100 ( .gnd(gnd), .vdd(vdd), .A(_3665_), .Y(_3666_) );
OAI21X1 OAI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_3488_), .B(_3486_), .C(_3477_), .Y(_3667_) );
NOR3X1 NOR3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3466_), .B(_2833_), .C(_3467_), .Y(_3668_) );
AOI21X1 AOI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_3471_), .B(_3468_), .C(_3668_), .Y(_3669_) );
INVX1 INVX1_452 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_19_), .Y(_3670_) );
INVX2 INVX2_101 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_3_), .Y(_3671_) );
NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_3671_), .B(_3459_), .Y(_3672_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_3459_), .B(_3671_), .Y(_3673_) );
OAI21X1 OAI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_3673_), .B(_3672_), .C(_3670_), .Y(_3674_) );
NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_3672_), .B(_3673_), .Y(_3675_) );
NAND2X1 NAND2X1_494 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_19_), .B(_3675_), .Y(_3676_) );
AOI21X1 AOI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_3674_), .B(_3676_), .C(_3464_), .Y(_3677_) );
INVX1 INVX1_453 ( .gnd(gnd), .vdd(vdd), .A(_3672_), .Y(_3678_) );
NAND2X1 NAND2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_3671_), .B(_3459_), .Y(_3679_) );
AOI21X1 AOI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_3679_), .B(_3678_), .C(module_0_W_19_), .Y(_3680_) );
NOR3X1 NOR3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_3672_), .B(_3670_), .C(_3673_), .Y(_3681_) );
NOR3X1 NOR3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_3467_), .B(_3681_), .C(_3680_), .Y(_3682_) );
OAI21X1 OAI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_3677_), .B(_3682_), .C(_3669_), .Y(_3683_) );
NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .B(_3677_), .Y(_3684_) );
OAI21X1 OAI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_3470_), .B(_3668_), .C(_3684_), .Y(_3685_) );
AOI21X1 AOI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_3683_), .B(_3685_), .C(bloque_datos_3_bF_buf3_), .Y(_3686_) );
INVX1 INVX1_454 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf2_), .Y(_3687_) );
INVX1 INVX1_455 ( .gnd(gnd), .vdd(vdd), .A(_3683_), .Y(_3688_) );
AOI21X1 AOI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_3464_), .B(_3462_), .C(_2790_), .Y(_3689_) );
OAI21X1 OAI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_3689_), .B(_2844_), .C(_3465_), .Y(_3690_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_3684_), .B(_3690_), .Y(_3691_) );
NOR3X1 NOR3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_3688_), .B(_3687_), .C(_3691_), .Y(_3692_) );
OAI21X1 OAI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_3692_), .B(_3686_), .C(_3479_), .Y(_3693_) );
OAI21X1 OAI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_3691_), .B(_3688_), .C(_3687_), .Y(_3694_) );
NAND3X1 NAND3X1_820 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf1_), .B(_3683_), .C(_3685_), .Y(_3695_) );
NAND3X1 NAND3X1_821 ( .gnd(gnd), .vdd(vdd), .A(_3476_), .B(_3695_), .C(_3694_), .Y(_3696_) );
AOI21X1 AOI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_3696_), .B(_3693_), .C(_3667_), .Y(_3697_) );
INVX2 INVX2_102 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .Y(_3698_) );
NAND3X1 NAND3X1_822 ( .gnd(gnd), .vdd(vdd), .A(_3667_), .B(_3696_), .C(_3693_), .Y(_3699_) );
AOI21X1 AOI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(_3698_), .C(bloque_datos_19_bF_buf3_), .Y(_3700_) );
INVX1 INVX1_456 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf2_), .Y(_3701_) );
INVX2 INVX2_103 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .Y(_3702_) );
NOR3X1 NOR3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_3701_), .B(_3697_), .C(_3702_), .Y(_3703_) );
OAI21X1 OAI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_3703_), .B(_3700_), .C(_3490_), .Y(_3704_) );
OAI21X1 OAI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_3702_), .B(_3697_), .C(_3701_), .Y(_3705_) );
NAND3X1 NAND3X1_823 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf1_), .B(_3699_), .C(_3698_), .Y(_3706_) );
NAND3X1 NAND3X1_824 ( .gnd(gnd), .vdd(vdd), .A(_3494_), .B(_3705_), .C(_3706_), .Y(_3707_) );
AOI21X1 AOI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_3707_), .B(_3704_), .C(_3666_), .Y(_3708_) );
NAND2X1 NAND2X1_496 ( .gnd(gnd), .vdd(vdd), .A(_3707_), .B(_3704_), .Y(_3709_) );
NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_3665_), .B(_3709_), .Y(_3710_) );
OAI21X1 OAI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_3710_), .B(_3708_), .C(bloque_datos_35_bF_buf4_), .Y(_3711_) );
INVX1 INVX1_457 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf3_), .Y(_3712_) );
INVX1 INVX1_458 ( .gnd(gnd), .vdd(vdd), .A(_3704_), .Y(_3713_) );
INVX1 INVX1_459 ( .gnd(gnd), .vdd(vdd), .A(_3707_), .Y(_3714_) );
OAI21X1 OAI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_3713_), .B(_3714_), .C(_3665_), .Y(_3715_) );
NAND3X1 NAND3X1_825 ( .gnd(gnd), .vdd(vdd), .A(_3707_), .B(_3704_), .C(_3666_), .Y(_3716_) );
NAND3X1 NAND3X1_826 ( .gnd(gnd), .vdd(vdd), .A(_3712_), .B(_3716_), .C(_3715_), .Y(_3717_) );
NAND3X1 NAND3X1_827 ( .gnd(gnd), .vdd(vdd), .A(_3506_), .B(_3717_), .C(_3711_), .Y(_3718_) );
OAI21X1 OAI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_3710_), .B(_3708_), .C(_3712_), .Y(_3719_) );
NAND3X1 NAND3X1_828 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf2_), .B(_3716_), .C(_3715_), .Y(_3720_) );
NAND3X1 NAND3X1_829 ( .gnd(gnd), .vdd(vdd), .A(_3503_), .B(_3720_), .C(_3719_), .Y(_3721_) );
NAND2X1 NAND2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_3718_), .B(_3721_), .Y(_3722_) );
NAND2X1 NAND2X1_498 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .B(_3664_), .Y(_3723_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_3664_), .B(_3722_), .Y(_3724_) );
NAND2X1 NAND2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_3723_), .B(_3724_), .Y(_3725_) );
XNOR2X1 XNOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_3725_), .B(bloque_datos_51_bF_buf4_), .Y(_3726_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_3726_), .B(_3663_), .Y(_3727_) );
NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_3509_), .B(_3513_), .Y(_3728_) );
INVX2 INVX2_104 ( .gnd(gnd), .vdd(vdd), .A(_3728_), .Y(_3729_) );
OAI21X1 OAI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_3512_), .B(_3729_), .C(_3726_), .Y(_3730_) );
AOI21X1 AOI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .B(_3727_), .C(_3662_), .Y(_3731_) );
INVX2 INVX2_105 ( .gnd(gnd), .vdd(vdd), .A(_3662_), .Y(_3732_) );
NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_3663_), .B(_3726_), .Y(_3733_) );
NAND2X1 NAND2X1_500 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf3_), .B(_3725_), .Y(_3734_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_3725_), .B(bloque_datos_51_bF_buf2_), .Y(_3735_) );
AOI21X1 AOI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_3734_), .B(_3735_), .C(_3514_), .Y(_3736_) );
NOR3X1 NOR3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_3732_), .B(_3736_), .C(_3733_), .Y(_3737_) );
OAI21X1 OAI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_3731_), .B(_3737_), .C(bloque_datos_67_bF_buf4_), .Y(_3738_) );
INVX1 INVX1_460 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf3_), .Y(_3739_) );
NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_3737_), .B(_3731_), .Y(_3740_) );
NAND2X1 NAND2X1_501 ( .gnd(gnd), .vdd(vdd), .A(_3739_), .B(_3740_), .Y(_3741_) );
NAND3X1 NAND3X1_830 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(_3738_), .C(_3741_), .Y(_3742_) );
OAI21X1 OAI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_3731_), .B(_3737_), .C(_3739_), .Y(_3743_) );
NAND2X1 NAND2X1_502 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf2_), .B(_3740_), .Y(_3744_) );
NAND3X1 NAND3X1_831 ( .gnd(gnd), .vdd(vdd), .A(_3526_), .B(_3743_), .C(_3744_), .Y(_3745_) );
AOI21X1 AOI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_3745_), .B(_3742_), .C(_3661_), .Y(_3746_) );
NAND3X1 NAND3X1_832 ( .gnd(gnd), .vdd(vdd), .A(_3661_), .B(_3745_), .C(_3742_), .Y(_3747_) );
INVX2 INVX2_106 ( .gnd(gnd), .vdd(vdd), .A(_3747_), .Y(_3748_) );
OAI21X1 OAI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .B(_3746_), .C(bloque_datos_83_bF_buf5_), .Y(_3749_) );
INVX1 INVX1_461 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf4_), .Y(_3750_) );
INVX2 INVX2_107 ( .gnd(gnd), .vdd(vdd), .A(_3746_), .Y(_3751_) );
NAND3X1 NAND3X1_833 ( .gnd(gnd), .vdd(vdd), .A(_3750_), .B(_3747_), .C(_3751_), .Y(_3752_) );
NAND3X1 NAND3X1_834 ( .gnd(gnd), .vdd(vdd), .A(_3541_), .B(_3752_), .C(_3749_), .Y(_3753_) );
INVX1 INVX1_462 ( .gnd(gnd), .vdd(vdd), .A(_3541_), .Y(_3754_) );
OAI21X1 OAI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .B(_3746_), .C(_3750_), .Y(_3755_) );
NAND3X1 NAND3X1_835 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf3_), .B(_3747_), .C(_3751_), .Y(_3756_) );
NAND3X1 NAND3X1_836 ( .gnd(gnd), .vdd(vdd), .A(_3754_), .B(_3756_), .C(_3755_), .Y(_3757_) );
AOI21X1 AOI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_3753_), .B(_3757_), .C(_3660_), .Y(_3758_) );
NAND3X1 NAND3X1_837 ( .gnd(gnd), .vdd(vdd), .A(_3660_), .B(_3753_), .C(_3757_), .Y(_3759_) );
INVX2 INVX2_108 ( .gnd(gnd), .vdd(vdd), .A(_3759_), .Y(_3760_) );
OAI21X1 OAI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_3760_), .B(_3758_), .C(_3659_), .Y(_3761_) );
INVX1 INVX1_463 ( .gnd(gnd), .vdd(vdd), .A(_3758_), .Y(_3762_) );
NAND3X1 NAND3X1_838 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_131_), .B(_3759_), .C(_3762_), .Y(_3763_) );
NAND2X1 NAND2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_3763_), .B(_3761_), .Y(_3764_) );
NAND2X1 NAND2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .B(_3764_), .Y(_3765_) );
INVX1 INVX1_464 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .Y(_3766_) );
NAND3X1 NAND3X1_839 ( .gnd(gnd), .vdd(vdd), .A(_3766_), .B(_3763_), .C(_3761_), .Y(_3767_) );
NAND3X1 NAND3X1_840 ( .gnd(gnd), .vdd(vdd), .A(_3767_), .B(_3765_), .C(_3658_), .Y(_3768_) );
INVX1 INVX1_465 ( .gnd(gnd), .vdd(vdd), .A(_3768_), .Y(_3769_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_3765_), .B(_3767_), .Y(_3770_) );
NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .B(_3770_), .Y(_3771_) );
OAI21X1 OAI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_3771_), .B(_3769_), .C(_3657_), .Y(_3772_) );
NOR3X1 NOR3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_3657_), .B(_3769_), .C(_3771_), .Y(_3773_) );
INVX2 INVX2_109 ( .gnd(gnd), .vdd(vdd), .A(_3773_), .Y(_3774_) );
NAND3X1 NAND3X1_841 ( .gnd(gnd), .vdd(vdd), .A(_3565_), .B(_3772_), .C(_3774_), .Y(_3775_) );
INVX1 INVX1_466 ( .gnd(gnd), .vdd(vdd), .A(_3565_), .Y(_3776_) );
INVX1 INVX1_467 ( .gnd(gnd), .vdd(vdd), .A(_3772_), .Y(_3777_) );
OAI21X1 OAI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_3777_), .B(_3773_), .C(_3776_), .Y(_3778_) );
NAND3X1 NAND3X1_842 ( .gnd(gnd), .vdd(vdd), .A(_3778_), .B(_3656_), .C(_3775_), .Y(_3779_) );
INVX1 INVX1_468 ( .gnd(gnd), .vdd(vdd), .A(_3779_), .Y(_3780_) );
AOI21X1 AOI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_3778_), .B(_3775_), .C(_3656_), .Y(_3781_) );
OAI21X1 OAI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_3780_), .B(_3781_), .C(_3654_), .Y(_3782_) );
NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_3781_), .B(_3780_), .Y(_3783_) );
NAND2X1 NAND2X1_505 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_163_), .B(_3783_), .Y(_3784_) );
NAND2X1 NAND2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_3782_), .B(_3784_), .Y(_3785_) );
NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_3575_), .B(_3785_), .Y(_3786_) );
INVX2 INVX2_110 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .Y(_3787_) );
OAI21X1 OAI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_3447_), .B(_3787_), .C(_3785_), .Y(_3788_) );
INVX2 INVX2_111 ( .gnd(gnd), .vdd(vdd), .A(_3788_), .Y(_3789_) );
NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_3786_), .B(_3789_), .Y(_3790_) );
OAI21X1 OAI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_3581_), .B(_3653_), .C(_3790_), .Y(_3791_) );
AOI21X1 AOI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .B(_3579_), .C(_3653_), .Y(_3792_) );
OAI21X1 OAI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_3789_), .B(_3786_), .C(_3792_), .Y(_3793_) );
NAND2X1 NAND2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_3793_), .B(_3791_), .Y(_3794_) );
NAND2X1 NAND2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_3652_), .B(_3794_), .Y(_3795_) );
NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_3652_), .B(_3794_), .Y(_3796_) );
INVX2 INVX2_112 ( .gnd(gnd), .vdd(vdd), .A(_3796_), .Y(_3797_) );
NAND3X1 NAND3X1_843 ( .gnd(gnd), .vdd(vdd), .A(_3588_), .B(_3795_), .C(_3797_), .Y(_3798_) );
INVX1 INVX1_469 ( .gnd(gnd), .vdd(vdd), .A(_3795_), .Y(_3799_) );
OAI21X1 OAI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_3799_), .B(_3796_), .C(_3585_), .Y(_3800_) );
NAND2X1 NAND2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_3800_), .B(_3798_), .Y(_3801_) );
NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_3651_), .B(_3801_), .Y(_3802_) );
INVX1 INVX1_470 ( .gnd(gnd), .vdd(vdd), .A(_3798_), .Y(_3803_) );
INVX1 INVX1_471 ( .gnd(gnd), .vdd(vdd), .A(_3800_), .Y(_3804_) );
OAI21X1 OAI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_3803_), .B(_3804_), .C(_3651_), .Y(_3805_) );
INVX1 INVX1_472 ( .gnd(gnd), .vdd(vdd), .A(_3805_), .Y(_3806_) );
OAI21X1 OAI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_3806_), .B(_3802_), .C(_3650_), .Y(_3807_) );
NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_3802_), .B(_3806_), .Y(_3808_) );
NAND2X1 NAND2X1_510 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_195_), .B(_3808_), .Y(_3809_) );
NAND2X1 NAND2X1_511 ( .gnd(gnd), .vdd(vdd), .A(_3807_), .B(_3809_), .Y(_3810_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_3810_), .B(_3649_), .Y(_3811_) );
AOI21X1 AOI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_3807_), .B(_3809_), .C(_3595_), .Y(_3812_) );
INVX1 INVX1_473 ( .gnd(gnd), .vdd(vdd), .A(_3812_), .Y(_3813_) );
NAND2X1 NAND2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_3813_), .B(_3811_), .Y(_3814_) );
NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_3648_), .B(_3814_), .Y(_3815_) );
NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_3649_), .B(_3810_), .Y(_3816_) );
OAI21X1 OAI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_3816_), .B(_3812_), .C(_3648_), .Y(_3817_) );
INVX2 INVX2_113 ( .gnd(gnd), .vdd(vdd), .A(_3817_), .Y(_3818_) );
OAI21X1 OAI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(_3815_), .B(_3818_), .C(_3646_), .Y(_3819_) );
INVX1 INVX1_474 ( .gnd(gnd), .vdd(vdd), .A(_3819_), .Y(_3820_) );
NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_3812_), .B(_3816_), .Y(_3821_) );
OAI21X1 OAI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_3647_), .B(_3600_), .C(_3821_), .Y(_3822_) );
NAND2X1 NAND2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_3817_), .B(_3822_), .Y(_3823_) );
NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_3646_), .B(_3823_), .Y(_3824_) );
NOR3X1 NOR3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_3645_), .B(_3824_), .C(_3820_), .Y(_3825_) );
NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_3818_), .B(_3815_), .Y(_3826_) );
NAND2X1 NAND2X1_514 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_211_), .B(_3826_), .Y(_3827_) );
AOI21X1 AOI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_3819_), .B(_3827_), .C(_3605_), .Y(_3828_) );
NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_3828_), .B(_3825_), .Y(_3829_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_3829_), .B(_3644_), .Y(_3830_) );
INVX1 INVX1_475 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .Y(_3831_) );
OAI21X1 OAI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_3825_), .B(_3828_), .C(_3831_), .Y(_3832_) );
INVX2 INVX2_114 ( .gnd(gnd), .vdd(vdd), .A(_3832_), .Y(_3833_) );
OAI21X1 OAI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(_3830_), .B(_3833_), .C(_3643_), .Y(_3834_) );
NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_3833_), .B(_3830_), .Y(_3835_) );
NAND2X1 NAND2X1_515 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_227_), .B(_3835_), .Y(_3836_) );
NAND3X1 NAND3X1_844 ( .gnd(gnd), .vdd(vdd), .A(_3618_), .B(_3834_), .C(_3836_), .Y(_3837_) );
NAND2X1 NAND2X1_516 ( .gnd(gnd), .vdd(vdd), .A(_3834_), .B(_3836_), .Y(_3838_) );
NAND2X1 NAND2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_3616_), .B(_3838_), .Y(_3839_) );
NAND3X1 NAND3X1_845 ( .gnd(gnd), .vdd(vdd), .A(_3642_), .B(_3837_), .C(_3839_), .Y(_3840_) );
INVX2 INVX2_115 ( .gnd(gnd), .vdd(vdd), .A(_3840_), .Y(_3841_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_3620_), .B(_3617_), .Y(_3842_) );
INVX1 INVX1_476 ( .gnd(gnd), .vdd(vdd), .A(_3837_), .Y(_3843_) );
AOI21X1 AOI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_3834_), .B(_3836_), .C(_3618_), .Y(_3844_) );
OAI21X1 OAI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_3843_), .B(_3844_), .C(_3842_), .Y(_3845_) );
INVX2 INVX2_116 ( .gnd(gnd), .vdd(vdd), .A(_3845_), .Y(_3846_) );
OAI21X1 OAI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_3846_), .B(_3841_), .C(_3641_), .Y(_3847_) );
NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_3841_), .B(_3846_), .Y(_3848_) );
NAND2X1 NAND2X1_518 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_243_), .B(_3848_), .Y(_3849_) );
NAND2X1 NAND2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_3847_), .B(_3849_), .Y(_3850_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_3850_), .B(_3625_), .Y(_3851_) );
INVX2 INVX2_117 ( .gnd(gnd), .vdd(vdd), .A(_3624_), .Y(_3852_) );
OAI21X1 OAI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_3852_), .B(_3444_), .C(_3850_), .Y(_3853_) );
AOI21X1 AOI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(_3851_), .C(_3640_), .Y(_3854_) );
INVX1 INVX1_477 ( .gnd(gnd), .vdd(vdd), .A(_3640_), .Y(_3855_) );
NAND2X1 NAND2X1_520 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(_3851_), .Y(_3856_) );
NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_3855_), .B(_3856_), .Y(_3857_) );
NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_3854_), .B(_3857_), .Y(_3858_) );
INVX2 INVX2_118 ( .gnd(gnd), .vdd(vdd), .A(_3858_), .Y(module_0_H_15_) );
NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_240_), .B(_3630_), .Y(_3859_) );
OAI21X1 OAI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_3632_), .B(_3443_), .C(_3859_), .Y(_3860_) );
NAND2X1 NAND2X1_521 ( .gnd(gnd), .vdd(vdd), .A(_3860_), .B(_3634_), .Y(_3861_) );
INVX2 INVX2_119 ( .gnd(gnd), .vdd(vdd), .A(_3861_), .Y(module_0_H_13_) );
NAND2X1 NAND2X1_522 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_240_), .B(_3630_), .Y(_3862_) );
INVX1 INVX1_478 ( .gnd(gnd), .vdd(vdd), .A(_3862_), .Y(_3863_) );
NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_3859_), .B(_3863_), .Y(module_0_H_0_) );
INVX1 INVX1_479 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_0_), .Y(module_0_H_12_) );
INVX1 INVX1_480 ( .gnd(gnd), .vdd(vdd), .A(_3634_), .Y(_3864_) );
OAI21X1 OAI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_3859_), .B(_3863_), .C(module_0_H_13_), .Y(_3865_) );
INVX2 INVX2_120 ( .gnd(gnd), .vdd(vdd), .A(_3865_), .Y(_3866_) );
AOI21X1 AOI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_3864_), .B(_3862_), .C(_3866_), .Y(module_0_H_1_) );
NAND3X1 NAND3X1_846 ( .gnd(gnd), .vdd(vdd), .A(_3626_), .B(_3864_), .C(_3638_), .Y(_3867_) );
INVX1 INVX1_481 ( .gnd(gnd), .vdd(vdd), .A(_3626_), .Y(_3868_) );
OAI21X1 OAI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_3639_), .B(_3868_), .C(_3634_), .Y(_3869_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_3869_), .B(_3867_), .Y(module_0_H_14_) );
NAND2X1 NAND2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_3866_), .B(module_0_H_14_), .Y(_3870_) );
INVX1 INVX1_482 ( .gnd(gnd), .vdd(vdd), .A(_3870_), .Y(_3871_) );
NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_3866_), .B(module_0_H_14_), .Y(_3872_) );
NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_3872_), .B(_3871_), .Y(module_0_H_2_) );
NOR3X1 NOR3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_3870_), .B(_3854_), .C(_3857_), .Y(_3873_) );
NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_3858_), .Y(_3874_) );
NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_3873_), .B(_3874_), .Y(module_0_H_3_) );
AOI21X1 AOI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_3847_), .B(_3849_), .C(_3637_), .Y(_3875_) );
OAI21X1 OAI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(_3855_), .B(_3875_), .C(_3851_), .Y(_3876_) );
INVX1 INVX1_483 ( .gnd(gnd), .vdd(vdd), .A(_3849_), .Y(_3877_) );
AOI21X1 AOI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_3642_), .B(_3839_), .C(_3843_), .Y(_3878_) );
OAI21X1 OAI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_3820_), .B(_3824_), .C(_3645_), .Y(_3879_) );
AOI21X1 AOI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3879_), .C(_3825_), .Y(_3880_) );
INVX1 INVX1_484 ( .gnd(gnd), .vdd(vdd), .A(_3648_), .Y(_3881_) );
AOI21X1 AOI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_3881_), .B(_3813_), .C(_3816_), .Y(_3882_) );
NAND2X1 NAND2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_3586_), .B(_3590_), .Y(_3883_) );
AOI21X1 AOI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_3883_), .B(_3800_), .C(_3803_), .Y(_3884_) );
INVX1 INVX1_485 ( .gnd(gnd), .vdd(vdd), .A(_3786_), .Y(_3885_) );
OAI21X1 OAI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(_3789_), .B(_3792_), .C(_3885_), .Y(_3886_) );
INVX1 INVX1_486 ( .gnd(gnd), .vdd(vdd), .A(_3886_), .Y(_3887_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_3779_), .B(_3775_), .Y(_3888_) );
NAND2X1 NAND2X1_525 ( .gnd(gnd), .vdd(vdd), .A(_3765_), .B(_3768_), .Y(_3889_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_3759_), .B(_3753_), .Y(_3890_) );
INVX2 INVX2_121 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .Y(_3891_) );
AOI21X1 AOI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_3743_), .B(_3744_), .C(_3526_), .Y(_3892_) );
AOI21X1 AOI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_3661_), .B(_3745_), .C(_3892_), .Y(_3893_) );
INVX2 INVX2_122 ( .gnd(gnd), .vdd(vdd), .A(_3743_), .Y(_3894_) );
AOI21X1 AOI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_3662_), .B(_3730_), .C(_3733_), .Y(_3895_) );
INVX1 INVX1_487 ( .gnd(gnd), .vdd(vdd), .A(_3725_), .Y(_3896_) );
NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf1_), .B(_3896_), .Y(_3897_) );
NAND2X1 NAND2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_3504_), .B(_3508_), .Y(_3898_) );
INVX1 INVX1_488 ( .gnd(gnd), .vdd(vdd), .A(_3718_), .Y(_3899_) );
AOI21X1 AOI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_3721_), .B(_3898_), .C(_3899_), .Y(_3900_) );
INVX2 INVX2_123 ( .gnd(gnd), .vdd(vdd), .A(_3719_), .Y(_3901_) );
AOI21X1 AOI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_3707_), .B(_3666_), .C(_3713_), .Y(_3902_) );
AOI21X1 AOI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_3695_), .B(_3694_), .C(_3476_), .Y(_3903_) );
AOI21X1 AOI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_3696_), .B(_3667_), .C(_3903_), .Y(_3904_) );
OAI21X1 OAI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(_3680_), .B(_3681_), .C(_3467_), .Y(_3905_) );
OAI21X1 OAI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(_3669_), .B(_3682_), .C(_3905_), .Y(_3906_) );
INVX1 INVX1_489 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_4_), .Y(_3907_) );
OAI21X1 OAI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_3459_), .B(_3671_), .C(_3907_), .Y(_3908_) );
NAND2X1 NAND2X1_527 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_4_), .B(_3672_), .Y(_3909_) );
AOI21X1 AOI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_3908_), .B(_3909_), .C(_2702_), .Y(_3910_) );
INVX1 INVX1_490 ( .gnd(gnd), .vdd(vdd), .A(_3908_), .Y(_3911_) );
NOR3X1 NOR3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_3671_), .B(_3907_), .C(_3459_), .Y(_3912_) );
NOR3X1 NOR3X1_102 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_0_), .B(_3912_), .C(_3911_), .Y(_3913_) );
OAI21X1 OAI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_3913_), .B(_3910_), .C(module_0_W_20_), .Y(_3914_) );
INVX1 INVX1_491 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_20_), .Y(_3915_) );
OAI21X1 OAI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(_3911_), .B(_3912_), .C(module_0_W_0_), .Y(_3916_) );
NAND3X1 NAND3X1_847 ( .gnd(gnd), .vdd(vdd), .A(_2702_), .B(_3908_), .C(_3909_), .Y(_3917_) );
NAND3X1 NAND3X1_848 ( .gnd(gnd), .vdd(vdd), .A(_3915_), .B(_3917_), .C(_3916_), .Y(_3918_) );
NAND3X1 NAND3X1_849 ( .gnd(gnd), .vdd(vdd), .A(_3674_), .B(_3918_), .C(_3914_), .Y(_3919_) );
OAI21X1 OAI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_3913_), .B(_3910_), .C(_3915_), .Y(_3920_) );
NAND3X1 NAND3X1_850 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_20_), .B(_3917_), .C(_3916_), .Y(_3921_) );
NAND3X1 NAND3X1_851 ( .gnd(gnd), .vdd(vdd), .A(_3680_), .B(_3921_), .C(_3920_), .Y(_3922_) );
NAND3X1 NAND3X1_852 ( .gnd(gnd), .vdd(vdd), .A(_3919_), .B(_3922_), .C(_3906_), .Y(_3923_) );
NAND3X1 NAND3X1_853 ( .gnd(gnd), .vdd(vdd), .A(_3464_), .B(_3674_), .C(_3676_), .Y(_3924_) );
AOI21X1 AOI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_3924_), .B(_3690_), .C(_3677_), .Y(_3925_) );
NAND3X1 NAND3X1_854 ( .gnd(gnd), .vdd(vdd), .A(_3680_), .B(_3918_), .C(_3914_), .Y(_3926_) );
NAND3X1 NAND3X1_855 ( .gnd(gnd), .vdd(vdd), .A(_3674_), .B(_3921_), .C(_3920_), .Y(_3927_) );
NAND3X1 NAND3X1_856 ( .gnd(gnd), .vdd(vdd), .A(_3925_), .B(_3926_), .C(_3927_), .Y(_3928_) );
XNOR2X1 XNOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .B(module_0_W_8_), .Y(_3929_) );
INVX1 INVX1_492 ( .gnd(gnd), .vdd(vdd), .A(_3929_), .Y(_3930_) );
NAND3X1 NAND3X1_857 ( .gnd(gnd), .vdd(vdd), .A(_3930_), .B(_3928_), .C(_3923_), .Y(_3931_) );
AOI21X1 AOI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_3926_), .B(_3927_), .C(_3925_), .Y(_3932_) );
AOI21X1 AOI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_3919_), .B(_3922_), .C(_3906_), .Y(_3933_) );
OAI21X1 OAI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_3932_), .B(_3933_), .C(_3929_), .Y(_3934_) );
AOI21X1 AOI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_3931_), .B(_3934_), .C(bloque_datos_4_bF_buf3_), .Y(_3935_) );
INVX1 INVX1_493 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf2_), .Y(_3936_) );
NAND3X1 NAND3X1_858 ( .gnd(gnd), .vdd(vdd), .A(_3929_), .B(_3928_), .C(_3923_), .Y(_3937_) );
OAI21X1 OAI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_3932_), .B(_3933_), .C(_3930_), .Y(_3938_) );
AOI21X1 AOI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_3937_), .B(_3938_), .C(_3936_), .Y(_3939_) );
OAI21X1 OAI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_3939_), .C(_3686_), .Y(_3940_) );
NAND3X1 NAND3X1_859 ( .gnd(gnd), .vdd(vdd), .A(_3936_), .B(_3937_), .C(_3938_), .Y(_3941_) );
NAND3X1 NAND3X1_860 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf1_), .B(_3931_), .C(_3934_), .Y(_3942_) );
NAND3X1 NAND3X1_861 ( .gnd(gnd), .vdd(vdd), .A(_3694_), .B(_3941_), .C(_3942_), .Y(_3943_) );
NAND3X1 NAND3X1_862 ( .gnd(gnd), .vdd(vdd), .A(_3904_), .B(_3943_), .C(_3940_), .Y(_3944_) );
AOI21X1 AOI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_3480_), .B(_3455_), .C(_3487_), .Y(_3945_) );
NOR3X1 NOR3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_3479_), .B(_3686_), .C(_3692_), .Y(_3946_) );
OAI21X1 OAI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_3946_), .B(_3945_), .C(_3693_), .Y(_3947_) );
OAI21X1 OAI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_3939_), .C(_3694_), .Y(_3948_) );
NAND3X1 NAND3X1_863 ( .gnd(gnd), .vdd(vdd), .A(_3686_), .B(_3941_), .C(_3942_), .Y(_3949_) );
NAND3X1 NAND3X1_864 ( .gnd(gnd), .vdd(vdd), .A(_3949_), .B(_3948_), .C(_3947_), .Y(_3950_) );
NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_24_), .B(module_0_W_8_), .Y(_3951_) );
INVX1 INVX1_494 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .Y(_3952_) );
NAND2X1 NAND2X1_528 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_24_), .B(module_0_W_8_), .Y(_3953_) );
NAND2X1 NAND2X1_529 ( .gnd(gnd), .vdd(vdd), .A(_3953_), .B(_3952_), .Y(_3954_) );
XNOR2X1 XNOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_2026_), .B(_3954_), .Y(_3955_) );
NAND3X1 NAND3X1_865 ( .gnd(gnd), .vdd(vdd), .A(_3955_), .B(_3944_), .C(_3950_), .Y(_3956_) );
AOI21X1 AOI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_3949_), .B(_3948_), .C(_3947_), .Y(_3957_) );
AOI21X1 AOI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_3943_), .B(_3940_), .C(_3904_), .Y(_3958_) );
INVX1 INVX1_495 ( .gnd(gnd), .vdd(vdd), .A(_3955_), .Y(_3959_) );
OAI21X1 OAI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_3957_), .B(_3958_), .C(_3959_), .Y(_3960_) );
AOI21X1 AOI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_3956_), .B(_3960_), .C(bloque_datos_20_bF_buf3_), .Y(_3961_) );
INVX1 INVX1_496 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf2_), .Y(_3962_) );
OAI21X1 OAI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_3957_), .B(_3958_), .C(_3955_), .Y(_3963_) );
NAND3X1 NAND3X1_866 ( .gnd(gnd), .vdd(vdd), .A(_3959_), .B(_3944_), .C(_3950_), .Y(_3964_) );
AOI21X1 AOI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_3964_), .B(_3963_), .C(_3962_), .Y(_3965_) );
OAI21X1 OAI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_3961_), .B(_3965_), .C(_3700_), .Y(_3966_) );
NAND3X1 NAND3X1_867 ( .gnd(gnd), .vdd(vdd), .A(_3962_), .B(_3964_), .C(_3963_), .Y(_3967_) );
NAND3X1 NAND3X1_868 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf1_), .B(_3956_), .C(_3960_), .Y(_3968_) );
NAND3X1 NAND3X1_869 ( .gnd(gnd), .vdd(vdd), .A(_3705_), .B(_3967_), .C(_3968_), .Y(_3969_) );
NAND3X1 NAND3X1_870 ( .gnd(gnd), .vdd(vdd), .A(_3969_), .B(_3966_), .C(_3902_), .Y(_3970_) );
OAI21X1 OAI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_3714_), .B(_3665_), .C(_3704_), .Y(_3971_) );
OAI21X1 OAI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_3961_), .B(_3965_), .C(_3705_), .Y(_3972_) );
NAND3X1 NAND3X1_871 ( .gnd(gnd), .vdd(vdd), .A(_3700_), .B(_3967_), .C(_3968_), .Y(_3973_) );
NAND3X1 NAND3X1_872 ( .gnd(gnd), .vdd(vdd), .A(_3973_), .B(_3971_), .C(_3972_), .Y(_3974_) );
INVX1 INVX1_497 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .Y(_3975_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_3954_), .B(_3975_), .Y(_3976_) );
NAND2X1 NAND2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_3975_), .B(_3954_), .Y(_3977_) );
NAND2X1 NAND2X1_531 ( .gnd(gnd), .vdd(vdd), .A(_3977_), .B(_3976_), .Y(_3978_) );
INVX2 INVX2_124 ( .gnd(gnd), .vdd(vdd), .A(_3978_), .Y(_3979_) );
XNOR2X1 XNOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_2057_), .B(_3979_), .Y(_3980_) );
NAND3X1 NAND3X1_873 ( .gnd(gnd), .vdd(vdd), .A(_3980_), .B(_3974_), .C(_3970_), .Y(_3981_) );
AOI21X1 AOI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_3973_), .B(_3972_), .C(_3971_), .Y(_172_) );
AOI21X1 AOI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_3969_), .B(_3966_), .C(_3902_), .Y(_173_) );
INVX1 INVX1_498 ( .gnd(gnd), .vdd(vdd), .A(_3980_), .Y(_174_) );
OAI21X1 OAI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_173_), .C(_174_), .Y(_175_) );
AOI21X1 AOI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_3981_), .B(_175_), .C(bloque_datos_36_bF_buf3_), .Y(_176_) );
INVX1 INVX1_499 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf2_), .Y(_177_) );
NAND3X1 NAND3X1_874 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_3974_), .C(_3970_), .Y(_178_) );
OAI21X1 OAI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_173_), .C(_3980_), .Y(_179_) );
AOI21X1 AOI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_179_), .C(_177_), .Y(_180_) );
OAI21X1 OAI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_180_), .C(_3901_), .Y(_181_) );
NAND3X1 NAND3X1_875 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_178_), .C(_179_), .Y(_182_) );
NAND3X1 NAND3X1_876 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf1_), .B(_3981_), .C(_175_), .Y(_183_) );
NAND3X1 NAND3X1_877 ( .gnd(gnd), .vdd(vdd), .A(_3719_), .B(_182_), .C(_183_), .Y(_184_) );
NAND3X1 NAND3X1_878 ( .gnd(gnd), .vdd(vdd), .A(_3900_), .B(_184_), .C(_181_), .Y(_185_) );
OAI21X1 OAI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(_3664_), .B(_3722_), .C(_3718_), .Y(_186_) );
OAI21X1 OAI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_180_), .C(_3719_), .Y(_187_) );
NAND3X1 NAND3X1_879 ( .gnd(gnd), .vdd(vdd), .A(_3901_), .B(_182_), .C(_183_), .Y(_188_) );
NAND3X1 NAND3X1_880 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_188_), .C(_187_), .Y(_189_) );
NAND2X1 NAND2X1_532 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf3_), .B(_3978_), .Y(_190_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_3978_), .B(bloque_datos_24_bF_buf2_), .Y(_191_) );
NAND2X1 NAND2X1_533 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .Y(_192_) );
INVX2 INVX2_125 ( .gnd(gnd), .vdd(vdd), .A(_192_), .Y(_193_) );
XNOR2X1 XNOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_2087_), .B(_193_), .Y(_194_) );
NAND3X1 NAND3X1_881 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_185_), .C(_189_), .Y(_195_) );
AOI21X1 AOI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_187_), .C(_186_), .Y(_196_) );
AOI21X1 AOI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_181_), .C(_3900_), .Y(_197_) );
INVX1 INVX1_500 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(_198_) );
OAI21X1 OAI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_197_), .C(_198_), .Y(_199_) );
AOI21X1 AOI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_199_), .C(bloque_datos_52_bF_buf4_), .Y(_200_) );
INVX1 INVX1_501 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf3_), .Y(_201_) );
NAND3X1 NAND3X1_882 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_185_), .C(_189_), .Y(_202_) );
OAI21X1 OAI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_197_), .C(_194_), .Y(_203_) );
AOI21X1 AOI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_203_), .C(_201_), .Y(_204_) );
OAI21X1 OAI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_204_), .C(_3897_), .Y(_205_) );
INVX2 INVX2_126 ( .gnd(gnd), .vdd(vdd), .A(_3897_), .Y(_206_) );
NAND3X1 NAND3X1_883 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_202_), .C(_203_), .Y(_207_) );
NAND3X1 NAND3X1_884 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf2_), .B(_195_), .C(_199_), .Y(_208_) );
NAND3X1 NAND3X1_885 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_207_), .C(_208_), .Y(_209_) );
NAND3X1 NAND3X1_886 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_3895_), .C(_205_), .Y(_210_) );
OAI21X1 OAI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_3736_), .B(_3732_), .C(_3727_), .Y(_211_) );
OAI21X1 OAI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_204_), .C(_206_), .Y(_212_) );
NAND3X1 NAND3X1_887 ( .gnd(gnd), .vdd(vdd), .A(_3897_), .B(_207_), .C(_208_), .Y(_213_) );
NAND3X1 NAND3X1_888 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_212_), .C(_211_), .Y(_214_) );
NAND2X1 NAND2X1_534 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf3_), .B(_192_), .Y(_215_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(bloque_datos_40_bF_buf2_), .Y(_216_) );
NAND2X1 NAND2X1_535 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_216_), .Y(_217_) );
INVX2 INVX2_127 ( .gnd(gnd), .vdd(vdd), .A(_217_), .Y(_218_) );
XNOR2X1 XNOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_2120_), .B(_218_), .Y(_219_) );
NAND3X1 NAND3X1_889 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_210_), .C(_214_), .Y(_220_) );
AOI21X1 AOI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_212_), .C(_211_), .Y(_221_) );
AOI21X1 AOI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_205_), .C(_3895_), .Y(_222_) );
INVX1 INVX1_502 ( .gnd(gnd), .vdd(vdd), .A(_219_), .Y(_223_) );
OAI21X1 OAI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_222_), .C(_223_), .Y(_224_) );
AOI21X1 AOI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_224_), .C(bloque_datos_68_bF_buf3_), .Y(_225_) );
INVX1 INVX1_503 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf2_), .Y(_226_) );
NAND3X1 NAND3X1_890 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_210_), .C(_214_), .Y(_227_) );
OAI21X1 OAI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_222_), .C(_219_), .Y(_228_) );
AOI21X1 AOI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_228_), .C(_226_), .Y(_229_) );
OAI21X1 OAI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_229_), .C(_3894_), .Y(_230_) );
NAND3X1 NAND3X1_891 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_227_), .C(_228_), .Y(_231_) );
NAND3X1 NAND3X1_892 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf1_), .B(_220_), .C(_224_), .Y(_232_) );
NAND3X1 NAND3X1_893 ( .gnd(gnd), .vdd(vdd), .A(_3743_), .B(_231_), .C(_232_), .Y(_233_) );
NAND3X1 NAND3X1_894 ( .gnd(gnd), .vdd(vdd), .A(_3893_), .B(_233_), .C(_230_), .Y(_234_) );
INVX1 INVX1_504 ( .gnd(gnd), .vdd(vdd), .A(_3661_), .Y(_235_) );
AOI21X1 AOI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_3738_), .B(_3741_), .C(_3530_), .Y(_236_) );
OAI21X1 OAI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_235_), .C(_3742_), .Y(_237_) );
OAI21X1 OAI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_229_), .C(_3743_), .Y(_238_) );
NAND3X1 NAND3X1_895 ( .gnd(gnd), .vdd(vdd), .A(_3894_), .B(_231_), .C(_232_), .Y(_239_) );
NAND3X1 NAND3X1_896 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_239_), .C(_238_), .Y(_240_) );
NAND2X1 NAND2X1_536 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf3_), .B(_217_), .Y(_241_) );
OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(bloque_datos_56_bF_buf2_), .Y(_242_) );
NAND2X1 NAND2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_242_), .Y(_243_) );
INVX2 INVX2_128 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_244_) );
XNOR2X1 XNOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_2153_), .B(_244_), .Y(_245_) );
NAND3X1 NAND3X1_897 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_234_), .C(_240_), .Y(_246_) );
AOI21X1 AOI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_238_), .C(_237_), .Y(_247_) );
AOI21X1 AOI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_230_), .C(_3893_), .Y(_248_) );
INVX1 INVX1_505 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_249_) );
OAI21X1 OAI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_248_), .C(_249_), .Y(_250_) );
AOI21X1 AOI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_250_), .C(bloque_datos_84_bF_buf4_), .Y(_251_) );
INVX1 INVX1_506 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf3_), .Y(_252_) );
NAND3X1 NAND3X1_898 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_234_), .C(_240_), .Y(_253_) );
OAI21X1 OAI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_248_), .C(_245_), .Y(_254_) );
AOI21X1 AOI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(_254_), .C(_252_), .Y(_255_) );
OAI21X1 OAI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_255_), .C(_3891_), .Y(_256_) );
NAND3X1 NAND3X1_899 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_253_), .C(_254_), .Y(_257_) );
NAND3X1 NAND3X1_900 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf2_), .B(_246_), .C(_250_), .Y(_258_) );
NAND3X1 NAND3X1_901 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .B(_257_), .C(_258_), .Y(_259_) );
NAND3X1 NAND3X1_902 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_259_), .C(_3890_), .Y(_260_) );
NAND2X1 NAND2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_3753_), .B(_3759_), .Y(_261_) );
OAI21X1 OAI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_255_), .C(_3755_), .Y(_262_) );
NAND3X1 NAND3X1_903 ( .gnd(gnd), .vdd(vdd), .A(_3891_), .B(_257_), .C(_258_), .Y(_263_) );
NAND3X1 NAND3X1_904 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf4_), .B(_244_), .Y(_265_) );
NAND2X1 NAND2X1_539 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf3_), .B(_244_), .Y(_266_) );
INVX1 INVX1_507 ( .gnd(gnd), .vdd(vdd), .A(_266_), .Y(_267_) );
NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_267_), .Y(_268_) );
XOR2X1 XOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(_268_), .Y(_269_) );
NAND3X1 NAND3X1_905 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_264_), .C(_260_), .Y(_270_) );
AOI21X1 AOI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_262_), .C(_261_), .Y(_271_) );
AOI21X1 AOI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_256_), .C(_3890_), .Y(_272_) );
INVX1 INVX1_508 ( .gnd(gnd), .vdd(vdd), .A(_269_), .Y(_273_) );
OAI21X1 OAI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_272_), .C(_273_), .Y(_274_) );
AOI21X1 AOI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_274_), .C(module_0_W_132_), .Y(_275_) );
INVX1 INVX1_509 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_132_), .Y(_276_) );
NAND3X1 NAND3X1_906 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_264_), .C(_260_), .Y(_277_) );
OAI21X1 OAI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_272_), .C(_269_), .Y(_278_) );
AOI21X1 AOI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_278_), .C(_276_), .Y(_279_) );
OAI21X1 OAI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_279_), .C(_3761_), .Y(_280_) );
INVX2 INVX2_129 ( .gnd(gnd), .vdd(vdd), .A(_3761_), .Y(_281_) );
NAND3X1 NAND3X1_907 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_277_), .C(_278_), .Y(_282_) );
NAND3X1 NAND3X1_908 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_132_), .B(_270_), .C(_274_), .Y(_283_) );
NAND3X1 NAND3X1_909 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_282_), .C(_283_), .Y(_284_) );
AOI21X1 AOI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_280_), .C(_3889_), .Y(_285_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_3768_), .B(_3765_), .Y(_286_) );
OAI21X1 OAI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_279_), .C(_281_), .Y(_287_) );
NAND3X1 NAND3X1_910 ( .gnd(gnd), .vdd(vdd), .A(_3761_), .B(_282_), .C(_283_), .Y(_288_) );
AOI21X1 AOI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_287_), .C(_286_), .Y(_289_) );
NAND2X1 NAND2X1_540 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf3_), .B(_268_), .Y(_290_) );
OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(bloque_datos_88_bF_buf2_), .Y(_291_) );
NAND2X1 NAND2X1_541 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_291_), .Y(_292_) );
OAI21X1 OAI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_289_), .C(_292_), .Y(_293_) );
AOI21X1 AOI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_283_), .C(_281_), .Y(_294_) );
NOR3X1 NOR3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_3761_), .C(_279_), .Y(_295_) );
OAI21X1 OAI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_294_), .C(_286_), .Y(_296_) );
NAND3X1 NAND3X1_911 ( .gnd(gnd), .vdd(vdd), .A(_3889_), .B(_284_), .C(_280_), .Y(_297_) );
INVX2 INVX2_130 ( .gnd(gnd), .vdd(vdd), .A(_292_), .Y(_298_) );
NAND3X1 NAND3X1_912 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_298_), .C(_296_), .Y(_299_) );
NAND2X1 NAND2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_299_), .Y(_300_) );
NAND3X1 NAND3X1_913 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_148_), .B(_2219_), .C(_300_), .Y(_301_) );
INVX1 INVX1_510 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_148_), .Y(_302_) );
AOI21X1 AOI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_296_), .C(_292_), .Y(_303_) );
NAND2X1 NAND2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_296_), .Y(_304_) );
OAI21X1 OAI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_298_), .C(_2219_), .Y(_305_) );
OAI21X1 OAI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_303_), .C(_302_), .Y(_306_) );
AOI21X1 AOI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_306_), .C(_3774_), .Y(_307_) );
OAI21X1 OAI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_303_), .C(module_0_W_148_), .Y(_308_) );
NAND3X1 NAND3X1_914 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_2219_), .C(_300_), .Y(_309_) );
AOI21X1 AOI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_308_), .C(_3773_), .Y(_310_) );
OAI21X1 OAI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_307_), .C(_3888_), .Y(_311_) );
NAND2X1 NAND2X1_544 ( .gnd(gnd), .vdd(vdd), .A(_3775_), .B(_3779_), .Y(_312_) );
NAND3X1 NAND3X1_915 ( .gnd(gnd), .vdd(vdd), .A(_3773_), .B(_309_), .C(_308_), .Y(_313_) );
NAND3X1 NAND3X1_916 ( .gnd(gnd), .vdd(vdd), .A(_3774_), .B(_301_), .C(_306_), .Y(_314_) );
NAND3X1 NAND3X1_917 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_313_), .C(_314_), .Y(_315_) );
NAND2X1 NAND2X1_545 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_136_), .B(_292_), .Y(_316_) );
OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(module_0_W_136_), .Y(_317_) );
NAND2X1 NAND2X1_546 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_317_), .Y(_318_) );
NAND3X1 NAND3X1_918 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_318_), .C(_311_), .Y(_319_) );
NAND2X1 NAND2X1_547 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_311_), .Y(_320_) );
INVX2 INVX2_131 ( .gnd(gnd), .vdd(vdd), .A(_318_), .Y(_321_) );
AOI21X1 AOI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_320_), .C(_2504_), .Y(_322_) );
NAND3X1 NAND3X1_919 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_164_), .B(_319_), .C(_322_), .Y(_323_) );
INVX1 INVX1_511 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_164_), .Y(_324_) );
AOI21X1 AOI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_314_), .C(_312_), .Y(_325_) );
NAND3X1 NAND3X1_920 ( .gnd(gnd), .vdd(vdd), .A(_3773_), .B(_301_), .C(_306_), .Y(_326_) );
NAND3X1 NAND3X1_921 ( .gnd(gnd), .vdd(vdd), .A(_3774_), .B(_309_), .C(_308_), .Y(_327_) );
AOI21X1 AOI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_327_), .C(_3888_), .Y(_328_) );
OAI21X1 OAI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_328_), .C(_321_), .Y(_329_) );
NAND3X1 NAND3X1_922 ( .gnd(gnd), .vdd(vdd), .A(_2252_), .B(_319_), .C(_329_), .Y(_330_) );
NAND2X1 NAND2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_330_), .Y(_331_) );
AOI21X1 AOI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_323_), .C(_3784_), .Y(_332_) );
INVX1 INVX1_512 ( .gnd(gnd), .vdd(vdd), .A(_3784_), .Y(_333_) );
NAND2X1 NAND2X1_549 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_164_), .B(_330_), .Y(_334_) );
NAND3X1 NAND3X1_923 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_319_), .C(_322_), .Y(_335_) );
AOI21X1 AOI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_335_), .C(_333_), .Y(_336_) );
OAI21X1 OAI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_332_), .C(_3887_), .Y(_337_) );
NAND3X1 NAND3X1_924 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_334_), .C(_335_), .Y(_338_) );
NAND3X1 NAND3X1_925 ( .gnd(gnd), .vdd(vdd), .A(_3784_), .B(_331_), .C(_323_), .Y(_339_) );
NAND3X1 NAND3X1_926 ( .gnd(gnd), .vdd(vdd), .A(_3886_), .B(_338_), .C(_339_), .Y(_340_) );
NAND2X1 NAND2X1_550 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_152_), .B(_318_), .Y(_341_) );
OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(module_0_W_152_), .Y(_342_) );
NAND2X1 NAND2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_342_), .Y(_343_) );
NAND3X1 NAND3X1_927 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_343_), .C(_337_), .Y(_344_) );
AOI21X1 AOI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_337_), .C(_343_), .Y(_345_) );
NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .B(_345_), .Y(_346_) );
NAND3X1 NAND3X1_928 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_180_), .B(_344_), .C(_346_), .Y(_347_) );
INVX1 INVX1_513 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_180_), .Y(_348_) );
NAND2X1 NAND2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_2285_), .B(_344_), .Y(_349_) );
OAI21X1 OAI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_345_), .C(_348_), .Y(_350_) );
AOI21X1 AOI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_347_), .C(_3797_), .Y(_351_) );
OAI21X1 OAI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_345_), .C(module_0_W_180_), .Y(_352_) );
NAND3X1 NAND3X1_929 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_344_), .C(_346_), .Y(_353_) );
AOI21X1 AOI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_353_), .C(_3796_), .Y(_354_) );
OAI21X1 OAI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_351_), .C(_3884_), .Y(_355_) );
OAI21X1 OAI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_3804_), .B(_3651_), .C(_3798_), .Y(_356_) );
NAND3X1 NAND3X1_930 ( .gnd(gnd), .vdd(vdd), .A(_3796_), .B(_352_), .C(_353_), .Y(_357_) );
NAND3X1 NAND3X1_931 ( .gnd(gnd), .vdd(vdd), .A(_3797_), .B(_350_), .C(_347_), .Y(_358_) );
NAND3X1 NAND3X1_932 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_356_), .C(_358_), .Y(_359_) );
NAND2X1 NAND2X1_553 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_168_), .B(_343_), .Y(_360_) );
OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(module_0_W_168_), .Y(_361_) );
NAND2X1 NAND2X1_554 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_361_), .Y(_362_) );
NAND3X1 NAND3X1_933 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_362_), .C(_355_), .Y(_363_) );
NAND2X1 NAND2X1_555 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_355_), .Y(_364_) );
INVX2 INVX2_132 ( .gnd(gnd), .vdd(vdd), .A(_362_), .Y(_365_) );
AOI21X1 AOI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_364_), .C(_2449_), .Y(_366_) );
NAND3X1 NAND3X1_934 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_196_), .B(_363_), .C(_366_), .Y(_367_) );
INVX1 INVX1_514 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_196_), .Y(_368_) );
AOI21X1 AOI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_358_), .C(_356_), .Y(_369_) );
NOR3X1 NOR3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_3884_), .C(_354_), .Y(_370_) );
OAI21X1 OAI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_369_), .C(_365_), .Y(_371_) );
NAND3X1 NAND3X1_935 ( .gnd(gnd), .vdd(vdd), .A(_2318_), .B(_363_), .C(_371_), .Y(_372_) );
NAND2X1 NAND2X1_556 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_372_), .Y(_373_) );
AOI21X1 AOI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_373_), .C(_3809_), .Y(_374_) );
INVX1 INVX1_515 ( .gnd(gnd), .vdd(vdd), .A(_3802_), .Y(_375_) );
NAND2X1 NAND2X1_557 ( .gnd(gnd), .vdd(vdd), .A(_3805_), .B(_375_), .Y(_376_) );
NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_3650_), .B(_376_), .Y(_377_) );
NAND2X1 NAND2X1_558 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_196_), .B(_372_), .Y(_378_) );
NAND3X1 NAND3X1_936 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_363_), .C(_366_), .Y(_379_) );
AOI21X1 AOI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_378_), .C(_377_), .Y(_380_) );
OAI21X1 OAI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_380_), .C(_3882_), .Y(_381_) );
OAI21X1 OAI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_3812_), .B(_3648_), .C(_3811_), .Y(_382_) );
NAND3X1 NAND3X1_937 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_379_), .C(_378_), .Y(_383_) );
NAND3X1 NAND3X1_938 ( .gnd(gnd), .vdd(vdd), .A(_3809_), .B(_367_), .C(_373_), .Y(_384_) );
NAND3X1 NAND3X1_939 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_384_), .C(_382_), .Y(_385_) );
NAND2X1 NAND2X1_559 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_381_), .Y(_386_) );
NAND2X1 NAND2X1_560 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_184_), .B(_362_), .Y(_387_) );
OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(module_0_W_184_), .Y(_388_) );
NAND2X1 NAND2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_388_), .Y(_389_) );
INVX2 INVX2_133 ( .gnd(gnd), .vdd(vdd), .A(_389_), .Y(_390_) );
OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_390_), .Y(_391_) );
AOI21X1 AOI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_381_), .C(_389_), .Y(_392_) );
NOR2X1 NOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_2428_), .B(_392_), .Y(_393_) );
NAND3X1 NAND3X1_940 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_212_), .B(_391_), .C(_393_), .Y(_394_) );
INVX1 INVX1_516 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_212_), .Y(_395_) );
OAI21X1 OAI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_390_), .C(_2351_), .Y(_396_) );
OAI21X1 OAI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_392_), .C(_395_), .Y(_397_) );
AOI21X1 AOI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_394_), .C(_3827_), .Y(_398_) );
OAI21X1 OAI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_392_), .C(module_0_W_212_), .Y(_399_) );
NAND3X1 NAND3X1_941 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_391_), .C(_393_), .Y(_400_) );
AOI21X1 AOI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_400_), .C(_3824_), .Y(_401_) );
OAI21X1 OAI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_401_), .C(_3880_), .Y(_402_) );
NAND3X1 NAND3X1_942 ( .gnd(gnd), .vdd(vdd), .A(_3605_), .B(_3819_), .C(_3827_), .Y(_403_) );
OAI21X1 OAI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_3831_), .B(_3828_), .C(_403_), .Y(_404_) );
NAND3X1 NAND3X1_943 ( .gnd(gnd), .vdd(vdd), .A(_3824_), .B(_399_), .C(_400_), .Y(_405_) );
NAND3X1 NAND3X1_944 ( .gnd(gnd), .vdd(vdd), .A(_3827_), .B(_397_), .C(_394_), .Y(_406_) );
INVX1 INVX1_517 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_0_), .Y(_4162_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .Y(_4163_) );
NAND2X1 NAND2X1_562 ( .gnd(gnd), .vdd(vdd), .A(nonce_iniciales[0]), .B(_4163_), .Y(_3983_) );
OAI21X1 OAI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_4162_), .B(_4163_), .C(_3983_), .Y(_3982__0_) );
INVX1 INVX1_518 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_1_), .Y(_3984_) );
NAND2X1 NAND2X1_563 ( .gnd(gnd), .vdd(vdd), .A(nonce_iniciales[1]), .B(_4163_), .Y(_3985_) );
OAI21X1 OAI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_4163_), .B(_3984_), .C(_3985_), .Y(_3982__1_) );
NAND2X1 NAND2X1_564 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_5_), .B(module_0_W_4_), .Y(_3986_) );
NAND2X1 NAND2X1_565 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_7_), .B(module_0_W_6_), .Y(_3987_) );
NOR2X1 NOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_3986_), .B(_3987_), .Y(_3988_) );
NAND2X1 NAND2X1_566 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_25_), .B(module_0_W_24_), .Y(_3989_) );
NAND2X1 NAND2X1_567 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_27_), .B(module_0_W_26_), .Y(_3990_) );
NOR2X1 NOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .B(_3990_), .Y(_3991_) );
INVX1 INVX1_519 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_2_), .Y(_3992_) );
OAI21X1 OAI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_4162_), .B(_3984_), .C(_3992_), .Y(_3993_) );
NAND3X1 NAND3X1_945 ( .gnd(gnd), .vdd(vdd), .A(_3993_), .B(_3988_), .C(_3991_), .Y(_3994_) );
INVX1 INVX1_520 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_29_), .Y(_3995_) );
INVX1 INVX1_521 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_28_), .Y(_3996_) );
NOR2X1 NOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_3995_), .B(_3996_), .Y(_3997_) );
INVX1 INVX1_522 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_31_), .Y(_3998_) );
INVX1 INVX1_523 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_30_), .Y(_3999_) );
NOR2X1 NOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_3998_), .B(_3999_), .Y(_4000_) );
NAND3X1 NAND3X1_946 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_3_), .B(_3997_), .C(_4000_), .Y(_4001_) );
NOR2X1 NOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_4001_), .B(_3994_), .Y(_4002_) );
NAND2X1 NAND2X1_568 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_17_), .B(module_0_W_16_), .Y(_4003_) );
NAND2X1 NAND2X1_569 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_19_), .B(module_0_W_18_), .Y(_4004_) );
NOR2X1 NOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_4003_), .B(_4004_), .Y(_4005_) );
NAND2X1 NAND2X1_570 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_22_), .B(module_0_W_21_), .Y(_4006_) );
NAND2X1 NAND2X1_571 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_23_), .B(module_0_W_20_), .Y(_4007_) );
NOR2X1 NOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_4006_), .B(_4007_), .Y(_4008_) );
NAND2X1 NAND2X1_572 ( .gnd(gnd), .vdd(vdd), .A(_4005_), .B(_4008_), .Y(_4009_) );
NAND2X1 NAND2X1_573 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_9_), .B(module_0_W_8_), .Y(_4010_) );
NAND2X1 NAND2X1_574 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_11_), .B(module_0_W_10_), .Y(_4011_) );
NOR2X1 NOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .B(_4011_), .Y(_4012_) );
NAND2X1 NAND2X1_575 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_15_), .B(module_0_W_14_), .Y(_4013_) );
NAND2X1 NAND2X1_576 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_13_), .B(module_0_W_12_), .Y(_4014_) );
NOR2X1 NOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_4013_), .B(_4014_), .Y(_4015_) );
NAND2X1 NAND2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_4012_), .B(_4015_), .Y(_4016_) );
NOR2X1 NOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4016_), .Y(_4017_) );
AOI21X1 AOI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_4017_), .B(_4002_), .C(_4163_), .Y(_4018_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_2_), .B(nonce_iniciales[2]), .S(inicio_bF_buf5), .Y(_4019_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_2_), .B(_4019_), .S(_4018__bF_buf1), .Y(_3982__2_) );
NAND2X1 NAND2X1_578 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_2_), .B(module_0_W_3_), .Y(_4020_) );
INVX1 INVX1_524 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_3_), .Y(_4021_) );
NAND2X1 NAND2X1_579 ( .gnd(gnd), .vdd(vdd), .A(_3992_), .B(_4021_), .Y(_4022_) );
NAND2X1 NAND2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_4020_), .B(_4022_), .Y(_4023_) );
NOR2X1 NOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf5), .B(nonce_iniciales[3]), .Y(_4024_) );
AOI21X1 AOI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_4023_), .B(_4018__bF_buf0), .C(_4024_), .Y(_3982__3_) );
XOR2X1 XOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_4020_), .B(module_0_W_4_), .Y(_4025_) );
NOR2X1 NOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf5), .B(nonce_iniciales[4]), .Y(_4026_) );
AOI21X1 AOI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_4025_), .B(_4018__bF_buf1), .C(_4026_), .Y(_3982__4_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_2_), .B(module_0_W_3_), .Y(_4027_) );
NAND2X1 NAND2X1_581 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_4_), .B(_4027_), .Y(_4028_) );
XOR2X1 XOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_4028_), .B(module_0_W_5_), .Y(_4029_) );
NOR2X1 NOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf5), .B(nonce_iniciales[5]), .Y(_4030_) );
AOI21X1 AOI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_4029_), .B(_4018__bF_buf0), .C(_4030_), .Y(_3982__5_) );
NOR2X1 NOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_3986_), .B(_4020_), .Y(_4031_) );
XNOR2X1 XNOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_4031_), .B(module_0_W_6_), .Y(_4032_) );
NOR2X1 NOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf5), .B(nonce_iniciales[6]), .Y(_4033_) );
AOI21X1 AOI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_4032_), .B(_4018__bF_buf1), .C(_4033_), .Y(_3982__6_) );
NOR2X1 NOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf5), .B(nonce_iniciales[7]), .Y(_4034_) );
NAND2X1 NAND2X1_582 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_6_), .B(_4031_), .Y(_4035_) );
XOR2X1 XOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_4035_), .B(module_0_W_7_), .Y(_4036_) );
AOI21X1 AOI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .B(_4018__bF_buf1), .C(_4034_), .Y(_3982__7_) );
NOR3X1 NOR3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_3986_), .B(_3987_), .C(_4020_), .Y(_4037_) );
XNOR2X1 XNOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_4037_), .B(module_0_W_8_), .Y(_4038_) );
NOR2X1 NOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf5), .B(nonce_iniciales[8]), .Y(_4039_) );
AOI21X1 AOI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .B(_4018__bF_buf0), .C(_4039_), .Y(_3982__8_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_5_), .B(module_0_W_4_), .Y(_4040_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_7_), .B(module_0_W_6_), .Y(_4041_) );
NAND3X1 NAND3X1_947 ( .gnd(gnd), .vdd(vdd), .A(_4040_), .B(_4041_), .C(_4027_), .Y(_4042_) );
INVX1 INVX1_525 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_9_), .Y(_4043_) );
INVX1 INVX1_526 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_8_), .Y(_4044_) );
OAI21X1 OAI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_4042_), .B(_4044_), .C(_4043_), .Y(_4045_) );
OAI21X1 OAI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .B(_4042_), .C(_4045_), .Y(_4046_) );
NOR2X1 NOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .B(nonce_iniciales[9]), .Y(_4047_) );
AOI21X1 AOI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_4046_), .B(_4018__bF_buf3), .C(_4047_), .Y(_3982__9_) );
NOR2X1 NOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .B(_4042_), .Y(_4048_) );
XNOR2X1 XNOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_4048_), .B(module_0_W_10_), .Y(_4049_) );
NOR2X1 NOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .B(nonce_iniciales[10]), .Y(_4050_) );
AOI21X1 AOI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_4049_), .B(_4018__bF_buf3), .C(_4050_), .Y(_3982__10_) );
NOR2X1 NOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .B(nonce_iniciales[11]), .Y(_4051_) );
NAND2X1 NAND2X1_583 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_10_), .B(_4048_), .Y(_4052_) );
OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_4052_), .B(module_0_W_11_), .Y(_4053_) );
NAND2X1 NAND2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_4017_), .B(_4002_), .Y(_4054_) );
NAND2X1 NAND2X1_585 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .B(_4054_), .Y(_4055_) );
AOI21X1 AOI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_11_), .B(_4052_), .C(_4055_), .Y(_4056_) );
AOI21X1 AOI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_4053_), .B(_4056_), .C(_4051_), .Y(_3982__11_) );
INVX2 INVX2_134 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_12_), .Y(_4057_) );
NAND2X1 NAND2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_4012_), .B(_4037_), .Y(_4058_) );
XNOR2X1 XNOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(_4057_), .Y(_4059_) );
NOR2X1 NOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .B(nonce_iniciales[12]), .Y(_4060_) );
AOI21X1 AOI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_4059_), .B(_4018__bF_buf3), .C(_4060_), .Y(_3982__12_) );
NOR2X1 NOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf5), .B(nonce_iniciales[13]), .Y(_4061_) );
INVX1 INVX1_527 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_13_), .Y(_4062_) );
NAND3X1 NAND3X1_948 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_11_), .B(module_0_W_10_), .C(_4048_), .Y(_4063_) );
NOR2X1 NOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_4057_), .B(_4063_), .Y(_4064_) );
NAND2X1 NAND2X1_587 ( .gnd(gnd), .vdd(vdd), .A(_4062_), .B(_4064_), .Y(_4065_) );
OAI21X1 OAI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(_4057_), .C(module_0_W_13_), .Y(_4066_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_4018__bF_buf3), .B(_4066_), .Y(_4067_) );
AOI21X1 AOI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_4065_), .B(_4067_), .C(_4061_), .Y(_3982__13_) );
INVX2 INVX2_135 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_14_), .Y(_4068_) );
OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(_4014_), .Y(_4069_) );
XNOR2X1 XNOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_4069_), .B(_4068_), .Y(_4070_) );
NOR2X1 NOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf5), .B(nonce_iniciales[14]), .Y(_4071_) );
AOI21X1 AOI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_4018__bF_buf1), .B(_4070_), .C(_4071_), .Y(_3982__14_) );
NOR2X1 NOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .B(nonce_iniciales[15]), .Y(_4072_) );
INVX1 INVX1_528 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_15_), .Y(_4073_) );
NOR2X1 NOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_4014_), .B(_4063_), .Y(_4074_) );
NAND3X1 NAND3X1_949 ( .gnd(gnd), .vdd(vdd), .A(_4073_), .B(module_0_W_14_), .C(_4074_), .Y(_4075_) );
OAI21X1 OAI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_4069_), .B(_4068_), .C(module_0_W_15_), .Y(_4076_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_4076_), .B(_4018__bF_buf3), .Y(_4077_) );
AOI21X1 AOI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_4075_), .B(_4077_), .C(_4072_), .Y(_3982__15_) );
OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .B(_4011_), .Y(_4078_) );
OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_4013_), .B(_4014_), .Y(_4079_) );
NOR3X1 NOR3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_4079_), .B(_4078_), .C(_4042_), .Y(_4080_) );
NAND2X1 NAND2X1_588 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_16_), .B(_4080_), .Y(_4081_) );
INVX1 INVX1_529 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_16_), .Y(_4082_) );
OAI21X1 OAI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_4016_), .B(_4042_), .C(_4082_), .Y(_4083_) );
NAND2X1 NAND2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_4083_), .B(_4081_), .Y(_4084_) );
NOR2X1 NOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf3), .B(nonce_iniciales[16]), .Y(_4085_) );
AOI21X1 AOI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(_4018__bF_buf2), .B(_4084_), .C(_4085_), .Y(_3982__16_) );
NAND3X1 NAND3X1_950 ( .gnd(gnd), .vdd(vdd), .A(_4012_), .B(_4015_), .C(_4037_), .Y(_4086_) );
NOR2X1 NOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_4082_), .B(_4086_), .Y(_4087_) );
XNOR2X1 XNOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_4087_), .B(module_0_W_17_), .Y(_4088_) );
NOR2X1 NOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf5), .B(nonce_iniciales[17]), .Y(_4089_) );
AOI21X1 AOI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_4018__bF_buf0), .B(_4088_), .C(_4089_), .Y(_3982__17_) );
INVX1 INVX1_530 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_18_), .Y(_4090_) );
INVX1 INVX1_531 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_17_), .Y(_4091_) );
OAI21X1 OAI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_4081_), .B(_4091_), .C(_4090_), .Y(_4092_) );
NAND3X1 NAND3X1_951 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_18_), .B(module_0_W_17_), .C(_4087_), .Y(_4093_) );
NAND2X1 NAND2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_4093_), .B(_4092_), .Y(_4094_) );
NOR2X1 NOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf3), .B(nonce_iniciales[18]), .Y(_4095_) );
AOI21X1 AOI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_4018__bF_buf2), .B(_4094_), .C(_4095_), .Y(_3982__18_) );
NOR2X1 NOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf3), .B(nonce_iniciales[19]), .Y(_4096_) );
OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_4093_), .B(module_0_W_19_), .Y(_4097_) );
AOI21X1 AOI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_19_), .B(_4093_), .C(_4055_), .Y(_4098_) );
AOI21X1 AOI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_4097_), .B(_4098_), .C(_4096_), .Y(_3982__19_) );
INVX1 INVX1_532 ( .gnd(gnd), .vdd(vdd), .A(_4005_), .Y(_4099_) );
NOR2X1 NOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_4099_), .B(_4086_), .Y(_4100_) );
NAND2X1 NAND2X1_591 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_20_), .B(_4100_), .Y(_4101_) );
INVX2 INVX2_136 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_20_), .Y(_4102_) );
OAI21X1 OAI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_4086_), .B(_4099_), .C(_4102_), .Y(_4103_) );
NAND2X1 NAND2X1_592 ( .gnd(gnd), .vdd(vdd), .A(_4103_), .B(_4101_), .Y(_4104_) );
NOR2X1 NOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf3), .B(nonce_iniciales[20]), .Y(_4105_) );
AOI21X1 AOI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_4018__bF_buf2), .B(_4104_), .C(_4105_), .Y(_3982__20_) );
INVX1 INVX1_533 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_21_), .Y(_4106_) );
INVX1 INVX1_534 ( .gnd(gnd), .vdd(vdd), .A(_4054_), .Y(_4107_) );
NAND2X1 NAND2X1_593 ( .gnd(gnd), .vdd(vdd), .A(_4005_), .B(_4080_), .Y(_4108_) );
NOR2X1 NOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_4102_), .B(_4108_), .Y(_4109_) );
AOI21X1 AOI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_4106_), .B(_4109_), .C(_4107_), .Y(_4110_) );
AOI21X1 AOI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_21_), .B(_4101_), .C(_4163_), .Y(_4111_) );
NOR2X1 NOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .B(nonce_iniciales[21]), .Y(_4112_) );
AOI21X1 AOI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_4111_), .B(_4110_), .C(_4112_), .Y(_3982__21_) );
NOR2X1 NOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_4106_), .B(_4102_), .Y(_4113_) );
INVX1 INVX1_535 ( .gnd(gnd), .vdd(vdd), .A(_4113_), .Y(_4114_) );
OAI21X1 OAI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_4108_), .B(_4114_), .C(module_0_W_22_), .Y(_4115_) );
INVX1 INVX1_536 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_22_), .Y(_4116_) );
NAND3X1 NAND3X1_952 ( .gnd(gnd), .vdd(vdd), .A(_4116_), .B(_4113_), .C(_4100_), .Y(_4117_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_4115_), .B(_4117_), .Y(_4118_) );
NOR2X1 NOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .B(nonce_iniciales[22]), .Y(_4119_) );
AOI21X1 AOI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_4018__bF_buf2), .B(_4118_), .C(_4119_), .Y(_3982__22_) );
NOR2X1 NOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf3), .B(nonce_iniciales[23]), .Y(_4120_) );
INVX1 INVX1_537 ( .gnd(gnd), .vdd(vdd), .A(_4006_), .Y(_4121_) );
NAND3X1 NAND3X1_953 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_20_), .B(_4121_), .C(_4100_), .Y(_4122_) );
OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_4122_), .B(module_0_W_23_), .Y(_4123_) );
AOI21X1 AOI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_23_), .B(_4122_), .C(_4055_), .Y(_4124_) );
AOI21X1 AOI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_4123_), .B(_4124_), .C(_4120_), .Y(_3982__23_) );
NOR2X1 NOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4086_), .Y(_4125_) );
XNOR2X1 XNOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_4125_), .B(module_0_W_24_), .Y(_4126_) );
NOR2X1 NOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf3), .B(nonce_iniciales[24]), .Y(_4127_) );
AOI21X1 AOI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(_4018__bF_buf2), .B(_4126_), .C(_4127_), .Y(_3982__24_) );
INVX1 INVX1_538 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_25_), .Y(_4128_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_4125_), .B(module_0_W_24_), .Y(_4129_) );
AOI21X1 AOI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(_4128_), .B(_4129_), .C(_4107_), .Y(_4130_) );
NAND2X1 NAND2X1_594 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_24_), .B(_4125_), .Y(_4131_) );
AOI21X1 AOI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_25_), .B(_4131_), .C(_4163_), .Y(_4132_) );
NOR2X1 NOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf3), .B(nonce_iniciales[25]), .Y(_4133_) );
AOI21X1 AOI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_4132_), .B(_4130_), .C(_4133_), .Y(_3982__25_) );
NOR3X1 NOR3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .B(_4009_), .C(_4086_), .Y(_4134_) );
XNOR2X1 XNOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_4134_), .B(module_0_W_26_), .Y(_4135_) );
NOR2X1 NOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .B(nonce_iniciales[26]), .Y(_4136_) );
AOI21X1 AOI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_4018__bF_buf2), .B(_4135_), .C(_4136_), .Y(_3982__26_) );
NOR2X1 NOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf3), .B(nonce_iniciales[27]), .Y(_4137_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_26_), .B(module_0_W_25_), .Y(_4138_) );
NAND3X1 NAND3X1_954 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_24_), .B(_4138_), .C(_4125_), .Y(_4139_) );
OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_4139_), .B(module_0_W_27_), .Y(_4140_) );
AOI21X1 AOI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_27_), .B(_4139_), .C(_4055_), .Y(_4141_) );
AOI21X1 AOI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_4140_), .B(_4141_), .C(_4137_), .Y(_3982__27_) );
INVX1 INVX1_539 ( .gnd(gnd), .vdd(vdd), .A(_3991_), .Y(_4142_) );
NOR3X1 NOR3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_4142_), .B(_4009_), .C(_4086_), .Y(_4143_) );
NAND2X1 NAND2X1_595 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_28_), .B(_4143_), .Y(_4144_) );
INVX1 INVX1_540 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .Y(_4145_) );
NAND3X1 NAND3X1_955 ( .gnd(gnd), .vdd(vdd), .A(_3991_), .B(_4145_), .C(_4080_), .Y(_4146_) );
NAND2X1 NAND2X1_596 ( .gnd(gnd), .vdd(vdd), .A(_3996_), .B(_4146_), .Y(_4147_) );
NAND2X1 NAND2X1_597 ( .gnd(gnd), .vdd(vdd), .A(_4144_), .B(_4147_), .Y(_4148_) );
NOR2X1 NOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .B(nonce_iniciales[28]), .Y(_4149_) );
AOI21X1 AOI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_4018__bF_buf3), .B(_4148_), .C(_4149_), .Y(_3982__28_) );
NOR2X1 NOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf10), .B(nonce_iniciales[29]), .Y(_4150_) );
OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_4144_), .B(module_0_W_29_), .Y(_4151_) );
AOI21X1 AOI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_29_), .B(_4144_), .C(_4055_), .Y(_4152_) );
AOI21X1 AOI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_4151_), .B(_4152_), .C(_4150_), .Y(_3982__29_) );
NAND3X1 NAND3X1_956 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_30_), .B(_3997_), .C(_4143_), .Y(_4153_) );
INVX1 INVX1_541 ( .gnd(gnd), .vdd(vdd), .A(_3997_), .Y(_4154_) );
OAI21X1 OAI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_4146_), .B(_4154_), .C(_3999_), .Y(_4155_) );
NAND2X1 NAND2X1_598 ( .gnd(gnd), .vdd(vdd), .A(_4153_), .B(_4155_), .Y(_4156_) );
NOR2X1 NOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf5), .B(nonce_iniciales[30]), .Y(_4157_) );
AOI21X1 AOI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_4018__bF_buf0), .B(_4156_), .C(_4157_), .Y(_3982__30_) );
NOR2X1 NOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf5), .B(nonce_iniciales[31]), .Y(_4158_) );
NOR2X1 NOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_4154_), .B(_4146_), .Y(_4159_) );
NAND3X1 NAND3X1_957 ( .gnd(gnd), .vdd(vdd), .A(_3998_), .B(module_0_W_30_), .C(_4159_), .Y(_4160_) );
AOI21X1 AOI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_31_), .B(_4153_), .C(_4055_), .Y(_4161_) );
AOI21X1 AOI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_4160_), .B(_4161_), .C(_4158_), .Y(_3982__31_) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__0_), .Q(module_0_W_0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__1_), .Q(module_0_W_1_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__2_), .Q(module_0_W_2_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__3_), .Q(module_0_W_3_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__4_), .Q(module_0_W_4_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__5_), .Q(module_0_W_5_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__6_), .Q(module_0_W_6_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__7_), .Q(module_0_W_7_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__8_), .Q(module_0_W_8_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__9_), .Q(module_0_W_9_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__10_), .Q(module_0_W_10_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__11_), .Q(module_0_W_11_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__12_), .Q(module_0_W_12_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__13_), .Q(module_0_W_13_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__14_), .Q(module_0_W_14_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__15_), .Q(module_0_W_15_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_3982__16_), .Q(module_0_W_16_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__17_), .Q(module_0_W_17_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_3982__18_), .Q(module_0_W_18_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__19_), .Q(module_0_W_19_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__20_), .Q(module_0_W_20_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3982__21_), .Q(module_0_W_21_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__22_), .Q(module_0_W_22_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3982__23_), .Q(module_0_W_23_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__24_), .Q(module_0_W_24_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3982__25_), .Q(module_0_W_25_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3982__26_), .Q(module_0_W_26_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3982__27_), .Q(module_0_W_27_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3982__28_), .Q(module_0_W_28_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_3982__29_), .Q(module_0_W_29_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__30_), .Q(module_0_W_30_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3982__31_), .Q(module_0_W_31_) );
INVX1 INVX1_542 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_4201_) );
INVX1 INVX1_543 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .Y(_4202_) );
INVX1 INVX1_544 ( .gnd(gnd), .vdd(vdd), .A(target[0]), .Y(_4203_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_4202_), .B(gnd), .C(_4203_), .D(vdd), .Y(_4204_) );
OAI21X1 OAI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .B(_4201_), .C(_4204_), .Y(_4205_) );
XOR2X1 XOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(vdd), .Y(_4206_) );
INVX2 INVX2_137 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .Y(_4207_) );
INVX1 INVX1_545 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_4208_) );
NAND2X1 NAND2X1_599 ( .gnd(gnd), .vdd(vdd), .A(_4207_), .B(_4208_), .Y(_4209_) );
NAND2X1 NAND2X1_600 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(gnd), .Y(_4210_) );
AOI21X1 AOI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_4209_), .B(_4210_), .C(_4206_), .Y(_4211_) );
INVX1 INVX1_546 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .Y(_4212_) );
NAND2X1 NAND2X1_601 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_4212_), .Y(_4213_) );
NAND2X1 NAND2X1_602 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_4207_), .Y(_4214_) );
OAI21X1 OAI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_4206_), .B(_4214_), .C(_4213_), .Y(_4215_) );
AOI21X1 AOI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_4205_), .B(_4211_), .C(_4215_), .Y(_4216_) );
INVX1 INVX1_547 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_15_), .Y(_4217_) );
INVX1 INVX1_548 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_14_), .Y(_4218_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_4217_), .B(target[7]), .C(target[6]), .D(_4218_), .Y(_4219_) );
INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .Y(_4220_) );
INVX2 INVX2_138 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .Y(_4221_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_4220_), .B(module_0_H_15_), .C(_4221_), .D(module_0_H_14_), .Y(_4222_) );
NOR2X1 NOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_4219_), .B(_4222_), .Y(_4223_) );
INVX2 INVX2_139 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_13_), .Y(_4224_) );
INVX1 INVX1_549 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_12_), .Y(_4225_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_4224_), .B(target[5]), .C(target[4]), .D(_4225_), .Y(_4226_) );
INVX2 INVX2_140 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .Y(_4227_) );
INVX1 INVX1_550 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .Y(_4228_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_4227_), .B(module_0_H_13_), .C(_4228_), .D(module_0_H_12_), .Y(_4229_) );
NOR2X1 NOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_4226_), .B(_4229_), .Y(_4230_) );
NAND2X1 NAND2X1_603 ( .gnd(gnd), .vdd(vdd), .A(_4223_), .B(_4230_), .Y(_4231_) );
NAND2X1 NAND2X1_604 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .B(_4224_), .Y(_4232_) );
NAND3X1 NAND3X1_958 ( .gnd(gnd), .vdd(vdd), .A(_4226_), .B(_4232_), .C(_4223_), .Y(_4233_) );
OAI21X1 OAI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_4216_), .B(_4231_), .C(_4233_), .Y(_4234_) );
INVX1 INVX1_551 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_17_), .Y(_4235_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_4202_), .B(module_0_H_17_), .C(_4203_), .D(module_0_H_16_), .Y(_4236_) );
OAI21X1 OAI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .B(_4235_), .C(_4236_), .Y(_4237_) );
XOR2X1 XOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(module_0_H_19_), .Y(_4238_) );
INVX1 INVX1_552 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_18_), .Y(_4239_) );
NAND2X1 NAND2X1_605 ( .gnd(gnd), .vdd(vdd), .A(_4207_), .B(_4239_), .Y(_4240_) );
NAND2X1 NAND2X1_606 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(module_0_H_18_), .Y(_4241_) );
AOI21X1 AOI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_4240_), .B(_4241_), .C(_4238_), .Y(_4242_) );
NAND2X1 NAND2X1_607 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_19_), .B(_4212_), .Y(_4164_) );
NAND2X1 NAND2X1_608 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_18_), .B(_4207_), .Y(_4165_) );
OAI21X1 OAI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(_4238_), .B(_4165_), .C(_4164_), .Y(_4166_) );
AOI21X1 AOI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_4237_), .B(_4242_), .C(_4166_), .Y(_4167_) );
INVX1 INVX1_553 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_23_), .Y(_4168_) );
INVX1 INVX1_554 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_22_), .Y(_4169_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_4168_), .B(target[7]), .C(target[6]), .D(_4169_), .Y(_4170_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_4220_), .B(module_0_H_23_), .C(_4221_), .D(module_0_H_22_), .Y(_4171_) );
NOR2X1 NOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_4170_), .B(_4171_), .Y(_4172_) );
NAND2X1 NAND2X1_609 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_21_), .B(_4227_), .Y(_4173_) );
NAND2X1 NAND2X1_610 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_20_), .B(_4228_), .Y(_4174_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_4173_), .B(_4174_), .Y(_4175_) );
INVX1 INVX1_555 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_20_), .Y(_4176_) );
NOR2X1 NOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_21_), .B(_4227_), .Y(_4177_) );
AOI21X1 AOI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_4176_), .C(_4177_), .Y(_4178_) );
NAND3X1 NAND3X1_959 ( .gnd(gnd), .vdd(vdd), .A(_4175_), .B(_4178_), .C(_4172_), .Y(_4179_) );
AOI21X1 AOI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_4173_), .B(_4174_), .C(_4177_), .Y(_4180_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_4220_), .B(module_0_H_23_), .C(_4221_), .D(module_0_H_22_), .Y(_4181_) );
NOR2X1 NOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_23_), .B(_4220_), .Y(_4182_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_4220_), .B(module_0_H_15_), .C(_4221_), .D(module_0_H_14_), .Y(_4183_) );
NOR2X1 NOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_15_), .B(_4220_), .Y(_4184_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_4181_), .B(_4182_), .C(_4183_), .D(_4184_), .Y(_4185_) );
AOI21X1 AOI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_4172_), .B(_4180_), .C(_4185_), .Y(_4186_) );
OAI21X1 OAI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_4167_), .B(_4179_), .C(_4186_), .Y(_4187_) );
NOR2X1 NOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf2), .B(_4187__bF_buf2), .Y(module_0_comparador_target_hash_0_terminado) );
INVX1 INVX1_556 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_0_), .Y(_4188_) );
NOR3X1 NOR3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf0), .B(_4188_), .C(_4187__bF_buf4), .Y(bounty_0_) );
INVX1 INVX1_557 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_1_), .Y(_4189_) );
NOR3X1 NOR3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf3), .B(_4189_), .C(_4187__bF_buf1), .Y(bounty_1_) );
INVX1 INVX1_558 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_2_), .Y(_4190_) );
NOR3X1 NOR3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf3), .B(_4190_), .C(_4187__bF_buf1), .Y(bounty_2_) );
INVX1 INVX1_559 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_3_), .Y(_4191_) );
NOR3X1 NOR3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf3), .B(_4191_), .C(_4187__bF_buf1), .Y(bounty_3_) );
INVX1 INVX1_560 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_4_), .Y(_4192_) );
NOR3X1 NOR3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf0), .B(_4192_), .C(_4187__bF_buf4), .Y(bounty_4_) );
INVX1 INVX1_561 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_5_), .Y(_4193_) );
NOR3X1 NOR3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf2), .B(_4193_), .C(_4187__bF_buf2), .Y(bounty_5_) );
INVX1 INVX1_562 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_6_), .Y(_4194_) );
NOR3X1 NOR3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf4), .B(_4194_), .C(_4187__bF_buf0), .Y(bounty_6_) );
INVX1 INVX1_563 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_7_), .Y(_4195_) );
NOR3X1 NOR3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf4), .B(_4195_), .C(_4187__bF_buf0), .Y(bounty_7_) );
INVX1 INVX1_564 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_4196_) );
NOR3X1 NOR3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf1), .B(_4196_), .C(_4187__bF_buf3), .Y(bounty_8_) );
NOR3X1 NOR3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf2), .B(_4201_), .C(_4187__bF_buf2), .Y(bounty_9_) );
NOR3X1 NOR3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf1), .B(_4208_), .C(_4187__bF_buf3), .Y(bounty_10_) );
INVX1 INVX1_565 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_4197_) );
NOR3X1 NOR3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf1), .B(_4197_), .C(_4187__bF_buf3), .Y(bounty_11_) );
NOR3X1 NOR3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf3), .B(_4225_), .C(_4187__bF_buf1), .Y(bounty_12_) );
NOR3X1 NOR3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf0), .B(_4224_), .C(_4187__bF_buf4), .Y(bounty_13_) );
NOR3X1 NOR3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf3), .B(_4218_), .C(_4187__bF_buf1), .Y(bounty_14_) );
NOR3X1 NOR3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf4), .B(_4217_), .C(_4187__bF_buf0), .Y(bounty_15_) );
INVX1 INVX1_566 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_16_), .Y(_4198_) );
NOR3X1 NOR3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf2), .B(_4198_), .C(_4187__bF_buf2), .Y(bounty_16_) );
NOR3X1 NOR3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf2), .B(_4235_), .C(_4187__bF_buf2), .Y(bounty_17_) );
NOR3X1 NOR3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf1), .B(_4239_), .C(_4187__bF_buf3), .Y(bounty_18_) );
INVX1 INVX1_567 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_19_), .Y(_4199_) );
NOR3X1 NOR3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf1), .B(_4199_), .C(_4187__bF_buf3), .Y(bounty_19_) );
NOR3X1 NOR3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf4), .B(_4176_), .C(_4187__bF_buf0), .Y(bounty_20_) );
INVX1 INVX1_568 ( .gnd(gnd), .vdd(vdd), .A(module_0_H_21_), .Y(_4200_) );
NOR3X1 NOR3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf4), .B(_4200_), .C(_4187__bF_buf0), .Y(bounty_21_) );
NOR3X1 NOR3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf0), .B(_4169_), .C(_4187__bF_buf4), .Y(bounty_22_) );
NOR3X1 NOR3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_4234__bF_buf0), .B(_4168_), .C(_4187__bF_buf4), .Y(bounty_23_) );
INVX1 INVX1_569 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf1_), .Y(_4243_) );
AOI21X1 AOI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_24_), .B(_4243_), .C(bloque_datos_80_bF_buf2_), .Y(_4244_) );
OAI21X1 OAI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_24_), .B(_4243_), .C(_4244_), .Y(module_0_W_136_) );
INVX1 INVX1_570 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf2_), .Y(_4245_) );
AOI21X1 AOI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_25_), .B(_4245_), .C(bloque_datos_81_bF_buf2_), .Y(_4246_) );
OAI21X1 OAI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_25_), .B(_4245_), .C(_4246_), .Y(module_0_W_137_) );
INVX1 INVX1_571 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf1_), .Y(_4247_) );
AOI21X1 AOI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_26_), .B(_4247_), .C(bloque_datos_82_bF_buf2_), .Y(_4248_) );
OAI21X1 OAI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_26_), .B(_4247_), .C(_4248_), .Y(module_0_W_138_) );
INVX1 INVX1_572 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf1_), .Y(_4249_) );
AOI21X1 AOI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_27_), .B(_4249_), .C(bloque_datos_83_bF_buf2_), .Y(_4250_) );
OAI21X1 OAI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_27_), .B(_4249_), .C(_4250_), .Y(module_0_W_139_) );
INVX1 INVX1_573 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf0_), .Y(_4251_) );
AOI21X1 AOI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_28_), .B(_4251_), .C(bloque_datos_84_bF_buf1_), .Y(_4252_) );
OAI21X1 OAI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_28_), .B(_4251_), .C(_4252_), .Y(module_0_W_140_) );
INVX1 INVX1_574 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf0_), .Y(_4253_) );
AOI21X1 AOI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_29_), .B(_4253_), .C(bloque_datos_85_bF_buf1_), .Y(_4254_) );
OAI21X1 OAI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_29_), .B(_4253_), .C(_4254_), .Y(module_0_W_141_) );
INVX1 INVX1_575 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf0_), .Y(_4255_) );
AOI21X1 AOI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_30_), .B(_4255_), .C(bloque_datos_86_bF_buf1_), .Y(_4256_) );
OAI21X1 OAI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_30_), .B(_4255_), .C(_4256_), .Y(module_0_W_142_) );
INVX1 INVX1_576 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .Y(_4257_) );
AOI21X1 AOI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_31_), .B(_4257_), .C(bloque_datos_87_bF_buf1_), .Y(_4258_) );
OAI21X1 OAI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_31_), .B(_4257_), .C(_4258_), .Y(module_0_W_143_) );
INVX1 INVX1_577 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf2_), .Y(_4259_) );
OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_16_), .B(bloque_datos_24_bF_buf1_), .Y(_4260_) );
NAND2X1 NAND2X1_611 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_16_), .B(bloque_datos_24_bF_buf0_), .Y(_4261_) );
NAND2X1 NAND2X1_612 ( .gnd(gnd), .vdd(vdd), .A(_4261_), .B(_4260_), .Y(_4262_) );
NAND2X1 NAND2X1_613 ( .gnd(gnd), .vdd(vdd), .A(_4259_), .B(_4262_), .Y(module_0_W_128_) );
INVX1 INVX1_578 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf1_), .Y(_4263_) );
AOI21X1 AOI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_17_), .B(_4263_), .C(bloque_datos_73_bF_buf2_), .Y(_4264_) );
OAI21X1 OAI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_17_), .B(_4263_), .C(_4264_), .Y(module_0_W_129_) );
INVX1 INVX1_579 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf2_), .Y(_4265_) );
OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_18_), .B(bloque_datos_26_bF_buf2_), .Y(_4266_) );
NAND2X1 NAND2X1_614 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_18_), .B(bloque_datos_26_bF_buf1_), .Y(_4267_) );
NAND2X1 NAND2X1_615 ( .gnd(gnd), .vdd(vdd), .A(_4267_), .B(_4266_), .Y(_4268_) );
NAND2X1 NAND2X1_616 ( .gnd(gnd), .vdd(vdd), .A(_4265_), .B(_4268_), .Y(module_0_W_130_) );
INVX1 INVX1_580 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf1_), .Y(_4269_) );
OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_19_), .B(bloque_datos_27_bF_buf1_), .Y(_4270_) );
NAND2X1 NAND2X1_617 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_19_), .B(bloque_datos_27_bF_buf0_), .Y(_4271_) );
NAND2X1 NAND2X1_618 ( .gnd(gnd), .vdd(vdd), .A(_4271_), .B(_4270_), .Y(_4272_) );
NAND2X1 NAND2X1_619 ( .gnd(gnd), .vdd(vdd), .A(_4269_), .B(_4272_), .Y(module_0_W_131_) );
INVX2 INVX2_141 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf1_), .Y(_4273_) );
AOI21X1 AOI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_20_), .B(_4273_), .C(bloque_datos_76_bF_buf1_), .Y(_4274_) );
OAI21X1 OAI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_20_), .B(_4273_), .C(_4274_), .Y(module_0_W_132_) );
INVX2 INVX2_142 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf1_), .Y(_4275_) );
AOI21X1 AOI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_21_), .B(_4275_), .C(bloque_datos_77_bF_buf1_), .Y(_4276_) );
OAI21X1 OAI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_21_), .B(_4275_), .C(_4276_), .Y(module_0_W_133_) );
INVX2 INVX2_143 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf0_), .Y(_4277_) );
AOI21X1 AOI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_22_), .B(_4277_), .C(bloque_datos_78_bF_buf1_), .Y(_4278_) );
OAI21X1 OAI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_22_), .B(_4277_), .C(_4278_), .Y(module_0_W_134_) );
INVX1 INVX1_581 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf1_), .Y(_4279_) );
AOI21X1 AOI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_23_), .B(_4279_), .C(bloque_datos_79_bF_buf2_), .Y(_4280_) );
OAI21X1 OAI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_23_), .B(_4279_), .C(_4280_), .Y(module_0_W_135_) );
INVX1 INVX1_582 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(_4281_) );
INVX1 INVX1_583 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf1_), .Y(_4282_) );
OAI21X1 OAI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_4281_), .B(bloque_datos_40_bF_buf1_), .C(_4282_), .Y(_4283_) );
AOI21X1 AOI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_4281_), .B(bloque_datos_40_bF_buf0_), .C(_4283_), .Y(_4284_) );
INVX1 INVX1_584 ( .gnd(gnd), .vdd(vdd), .A(_4284_), .Y(module_0_W_144_) );
INVX1 INVX1_585 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(_4285_) );
INVX1 INVX1_586 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf2_), .Y(_4286_) );
OAI21X1 OAI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_4285_), .B(bloque_datos_41_bF_buf1_), .C(_4286_), .Y(_4287_) );
AOI21X1 AOI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_4285_), .B(bloque_datos_41_bF_buf0_), .C(_4287_), .Y(_4288_) );
INVX1 INVX1_587 ( .gnd(gnd), .vdd(vdd), .A(_4288_), .Y(module_0_W_145_) );
INVX1 INVX1_588 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf0_), .Y(_4289_) );
INVX1 INVX1_589 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf1_), .Y(_4290_) );
OAI21X1 OAI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_4289_), .B(bloque_datos_42_bF_buf1_), .C(_4290_), .Y(_4291_) );
AOI21X1 AOI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_4289_), .B(bloque_datos_42_bF_buf0_), .C(_4291_), .Y(_4292_) );
INVX1 INVX1_590 ( .gnd(gnd), .vdd(vdd), .A(_4292_), .Y(module_0_W_146_) );
INVX1 INVX1_591 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf0_), .Y(_4293_) );
INVX1 INVX1_592 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf0_), .Y(_4294_) );
OAI21X1 OAI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_4293_), .B(bloque_datos_43_bF_buf1_), .C(_4294_), .Y(_4295_) );
AOI21X1 AOI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(_4293_), .B(bloque_datos_43_bF_buf0_), .C(_4295_), .Y(_4296_) );
INVX1 INVX1_593 ( .gnd(gnd), .vdd(vdd), .A(_4296_), .Y(module_0_W_147_) );
INVX1 INVX1_594 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf0_), .Y(_4297_) );
INVX1 INVX1_595 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf0_), .Y(_4298_) );
OAI21X1 OAI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_4297_), .B(bloque_datos_44_bF_buf1_), .C(_4298_), .Y(_4299_) );
AOI21X1 AOI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_4297_), .B(bloque_datos_44_bF_buf0_), .C(_4299_), .Y(_4300_) );
INVX1 INVX1_596 ( .gnd(gnd), .vdd(vdd), .A(_4300_), .Y(module_0_W_148_) );
INVX1 INVX1_597 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf0_), .Y(_4301_) );
INVX1 INVX1_598 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf0_), .Y(_4302_) );
OAI21X1 OAI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_4301_), .B(bloque_datos_45_bF_buf1_), .C(_4302_), .Y(_4303_) );
AOI21X1 AOI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_4301_), .B(bloque_datos_45_bF_buf0_), .C(_4303_), .Y(_4304_) );
INVX1 INVX1_599 ( .gnd(gnd), .vdd(vdd), .A(_4304_), .Y(module_0_W_149_) );
INVX1 INVX1_600 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf0_), .Y(_4305_) );
INVX1 INVX1_601 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf0_), .Y(_4306_) );
OAI21X1 OAI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_4305_), .B(bloque_datos_46_bF_buf1_), .C(_4306_), .Y(_4307_) );
AOI21X1 AOI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_4305_), .B(bloque_datos_46_bF_buf0_), .C(_4307_), .Y(_4308_) );
INVX2 INVX2_144 ( .gnd(gnd), .vdd(vdd), .A(_4308_), .Y(module_0_W_150_) );
INVX1 INVX1_602 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[7]), .Y(_4309_) );
INVX1 INVX1_603 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf1_), .Y(_4310_) );
OAI21X1 OAI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_4309_), .B(bloque_datos_47_bF_buf2_), .C(_4310_), .Y(_4311_) );
AOI21X1 AOI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_4309_), .B(bloque_datos_47_bF_buf1_), .C(_4311_), .Y(_4312_) );
INVX2 INVX2_145 ( .gnd(gnd), .vdd(vdd), .A(_4312_), .Y(module_0_W_151_) );
AOI21X1 AOI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_4261_), .B(_4260_), .C(bloque_datos_72_bF_buf1_), .Y(_4313_) );
XNOR2X1 XNOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .B(bloque_datos_48_bF_buf1_), .Y(_4314_) );
NAND2X1 NAND2X1_620 ( .gnd(gnd), .vdd(vdd), .A(_4314_), .B(_4313_), .Y(module_0_W_152_) );
XOR2X1 XOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .B(bloque_datos_49_bF_buf2_), .Y(_4315_) );
NOR2X1 NOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_4315_), .B(module_0_W_129_), .Y(_4316_) );
INVX1 INVX1_604 ( .gnd(gnd), .vdd(vdd), .A(_4316_), .Y(module_0_W_153_) );
AOI21X1 AOI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_4267_), .B(_4266_), .C(bloque_datos_74_bF_buf1_), .Y(_4317_) );
XNOR2X1 XNOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .B(bloque_datos_50_bF_buf1_), .Y(_4318_) );
NAND2X1 NAND2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_4318_), .B(_4317_), .Y(module_0_W_154_) );
AOI21X1 AOI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_4271_), .B(_4270_), .C(bloque_datos_75_bF_buf0_), .Y(_4319_) );
XNOR2X1 XNOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .B(bloque_datos_51_bF_buf0_), .Y(_4320_) );
NAND2X1 NAND2X1_622 ( .gnd(gnd), .vdd(vdd), .A(_4320_), .B(_4319_), .Y(module_0_W_155_) );
INVX1 INVX1_605 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_20_), .Y(_4321_) );
INVX1 INVX1_606 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf0_), .Y(_4322_) );
OAI21X1 OAI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_4321_), .B(bloque_datos_28_bF_buf0_), .C(_4322_), .Y(_4323_) );
AOI21X1 AOI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_4321_), .B(bloque_datos_28_bF_buf4_), .C(_4323_), .Y(_4324_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf0_), .B(bloque_datos_52_bF_buf1_), .Y(_4325_) );
NOR2X1 NOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf3_), .B(bloque_datos_52_bF_buf0_), .Y(_4326_) );
OAI21X1 OAI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_4325_), .B(_4326_), .C(_4324_), .Y(module_0_W_156_) );
XOR2X1 XOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf0_), .B(bloque_datos_53_bF_buf0_), .Y(_4327_) );
NOR2X1 NOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_4327_), .B(module_0_W_133_), .Y(_4328_) );
INVX1 INVX1_607 ( .gnd(gnd), .vdd(vdd), .A(_4328_), .Y(module_0_W_157_) );
XOR2X1 XOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf0_), .B(bloque_datos_54_bF_buf0_), .Y(_4329_) );
NOR2X1 NOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_4329_), .B(module_0_W_134_), .Y(_4330_) );
INVX1 INVX1_608 ( .gnd(gnd), .vdd(vdd), .A(_4330_), .Y(module_0_W_158_) );
XOR2X1 XOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[15]), .B(bloque_datos[55]), .Y(_4331_) );
NOR2X1 NOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_4331_), .B(module_0_W_135_), .Y(_4332_) );
INVX1 INVX1_609 ( .gnd(gnd), .vdd(vdd), .A(_4332_), .Y(module_0_W_159_) );
XOR2X1 XOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_24_), .B(bloque_datos_32_bF_buf0_), .Y(_4333_) );
NOR2X1 NOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf1_), .B(_4333_), .Y(_4334_) );
XNOR2X1 XNOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf0_), .B(bloque_datos_56_bF_buf1_), .Y(_4335_) );
NAND2X1 NAND2X1_623 ( .gnd(gnd), .vdd(vdd), .A(_4335_), .B(_4334_), .Y(module_0_W_160_) );
INVX1 INVX1_610 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_25_), .Y(_4336_) );
INVX1 INVX1_611 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf1_), .Y(_4337_) );
OAI21X1 OAI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(_4336_), .B(bloque_datos_33_bF_buf1_), .C(_4337_), .Y(_4338_) );
AOI21X1 AOI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_4336_), .B(bloque_datos_33_bF_buf0_), .C(_4338_), .Y(_4339_) );
XNOR2X1 XNOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .B(bloque_datos_57_bF_buf1_), .Y(_4340_) );
NAND2X1 NAND2X1_624 ( .gnd(gnd), .vdd(vdd), .A(_4340_), .B(_4339_), .Y(module_0_W_161_) );
XOR2X1 XOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_26_), .B(bloque_datos_34_bF_buf0_), .Y(_4341_) );
NOR2X1 NOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf1_), .B(_4341_), .Y(_4342_) );
XNOR2X1 XNOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .B(bloque_datos_58_bF_buf1_), .Y(_4343_) );
NAND2X1 NAND2X1_625 ( .gnd(gnd), .vdd(vdd), .A(_4343_), .B(_4342_), .Y(module_0_W_162_) );
XOR2X1 XOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_27_), .B(bloque_datos_35_bF_buf0_), .Y(_4344_) );
NOR2X1 NOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf1_), .B(_4344_), .Y(_4345_) );
XNOR2X1 XNOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf0_), .B(bloque_datos_59_bF_buf1_), .Y(_4346_) );
NAND2X1 NAND2X1_626 ( .gnd(gnd), .vdd(vdd), .A(_4346_), .B(_4345_), .Y(module_0_W_163_) );
XOR2X1 XOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf0_), .B(bloque_datos_60_bF_buf0_), .Y(_4347_) );
NOR2X1 NOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_4347_), .B(module_0_W_140_), .Y(_4348_) );
INVX1 INVX1_612 ( .gnd(gnd), .vdd(vdd), .A(_4348_), .Y(module_0_W_164_) );
XOR2X1 XOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf0_), .B(bloque_datos_61_bF_buf1_), .Y(_4349_) );
NOR2X1 NOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_4349_), .B(module_0_W_141_), .Y(_4350_) );
INVX1 INVX1_613 ( .gnd(gnd), .vdd(vdd), .A(_4350_), .Y(module_0_W_165_) );
XOR2X1 XOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf0_), .B(bloque_datos_62_bF_buf0_), .Y(_4351_) );
NOR2X1 NOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_4351_), .B(module_0_W_142_), .Y(_4352_) );
INVX2 INVX2_146 ( .gnd(gnd), .vdd(vdd), .A(_4352_), .Y(module_0_W_166_) );
XOR2X1 XOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf0_), .B(bloque_datos[63]), .Y(_4353_) );
NOR2X1 NOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_4353_), .B(module_0_W_143_), .Y(_4354_) );
INVX1 INVX1_614 ( .gnd(gnd), .vdd(vdd), .A(_4354_), .Y(module_0_W_167_) );
XNOR2X1 XNOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf4_), .B(bloque_datos_64_bF_buf1_), .Y(_4355_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_4284_), .B(_4355_), .Y(_4356_) );
INVX2 INVX2_147 ( .gnd(gnd), .vdd(vdd), .A(_4356_), .Y(module_0_W_168_) );
XNOR2X1 XNOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf0_), .B(bloque_datos_65_bF_buf1_), .Y(_4357_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_4288_), .B(_4357_), .Y(_4358_) );
INVX1 INVX1_615 ( .gnd(gnd), .vdd(vdd), .A(_4358_), .Y(module_0_W_169_) );
XNOR2X1 XNOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf0_), .B(bloque_datos_66_bF_buf1_), .Y(_4359_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_4292_), .B(_4359_), .Y(_4360_) );
INVX1 INVX1_616 ( .gnd(gnd), .vdd(vdd), .A(_4360_), .Y(module_0_W_170_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf4_), .B(bloque_datos_67_bF_buf1_), .Y(_4361_) );
NOR2X1 NOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf3_), .B(bloque_datos_67_bF_buf0_), .Y(_4362_) );
OAI21X1 OAI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_4361_), .B(_4362_), .C(_4296_), .Y(module_0_W_171_) );
INVX2 INVX2_148 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf0_), .Y(_4363_) );
NOR2X1 NOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_4273_), .B(_4363_), .Y(_4364_) );
NOR2X1 NOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf3_), .B(bloque_datos_68_bF_buf3_), .Y(_4365_) );
OAI21X1 OAI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(_4364_), .B(_4365_), .C(_4300_), .Y(module_0_W_172_) );
INVX2 INVX2_149 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf0_), .Y(_4366_) );
NOR2X1 NOR2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_4275_), .B(_4366_), .Y(_4367_) );
NOR2X1 NOR2X1_340 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf0_), .B(bloque_datos_69_bF_buf3_), .Y(_4368_) );
OAI21X1 OAI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_4367_), .B(_4368_), .C(_4304_), .Y(module_0_W_173_) );
INVX2 INVX2_150 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf0_), .Y(_4369_) );
NOR2X1 NOR2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_4277_), .B(_4369_), .Y(_4370_) );
NOR2X1 NOR2X1_342 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf3_), .B(bloque_datos_70_bF_buf3_), .Y(_4371_) );
OAI21X1 OAI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_4370_), .B(_4371_), .C(_4308_), .Y(module_0_W_174_) );
XNOR2X1 XNOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf0_), .B(bloque_datos_71_bF_buf1_), .Y(_4372_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_4312_), .B(_4372_), .Y(_4373_) );
INVX1 INVX1_617 ( .gnd(gnd), .vdd(vdd), .A(_4373_), .Y(module_0_W_175_) );
XNOR2X1 XNOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf4_), .B(bloque_datos_72_bF_buf0_), .Y(_4374_) );
NAND3X1 NAND3X1_960 ( .gnd(gnd), .vdd(vdd), .A(_4314_), .B(_4374_), .C(_4313_), .Y(module_0_W_176_) );
INVX1 INVX1_618 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_17_), .Y(_4375_) );
NAND2X1 NAND2X1_627 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf3_), .B(_4375_), .Y(_4376_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_4264_), .B(_4376_), .Y(_4377_) );
INVX1 INVX1_619 ( .gnd(gnd), .vdd(vdd), .A(_4315_), .Y(_4378_) );
XNOR2X1 XNOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf3_), .B(bloque_datos_73_bF_buf1_), .Y(_4379_) );
NAND3X1 NAND3X1_961 ( .gnd(gnd), .vdd(vdd), .A(_4378_), .B(_4379_), .C(_4377_), .Y(module_0_W_177_) );
XNOR2X1 XNOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf4_), .B(bloque_datos_74_bF_buf0_), .Y(_4380_) );
NAND3X1 NAND3X1_962 ( .gnd(gnd), .vdd(vdd), .A(_4318_), .B(_4380_), .C(_4317_), .Y(module_0_W_178_) );
XNOR2X1 XNOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf4_), .B(bloque_datos_75_bF_buf4_), .Y(_4381_) );
NAND3X1 NAND3X1_963 ( .gnd(gnd), .vdd(vdd), .A(_4320_), .B(_4381_), .C(_4319_), .Y(module_0_W_179_) );
XOR2X1 XOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf3_), .B(bloque_datos_76_bF_buf4_), .Y(_4382_) );
NOR2X1 NOR2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_4382_), .B(module_0_W_156_), .Y(_4383_) );
INVX1 INVX1_620 ( .gnd(gnd), .vdd(vdd), .A(_4383_), .Y(module_0_W_180_) );
INVX1 INVX1_621 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_21_), .Y(_4384_) );
INVX1 INVX1_622 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf0_), .Y(_4385_) );
OAI21X1 OAI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_4384_), .B(bloque_datos_29_bF_buf4_), .C(_4385_), .Y(_4386_) );
AOI21X1 AOI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_4384_), .B(bloque_datos_29_bF_buf3_), .C(_4386_), .Y(_4387_) );
INVX1 INVX1_623 ( .gnd(gnd), .vdd(vdd), .A(_4327_), .Y(_4388_) );
XNOR2X1 XNOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf3_), .B(bloque_datos_77_bF_buf4_), .Y(_4389_) );
NAND3X1 NAND3X1_964 ( .gnd(gnd), .vdd(vdd), .A(_4388_), .B(_4389_), .C(_4387_), .Y(module_0_W_181_) );
XNOR2X1 XNOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf3_), .B(bloque_datos_78_bF_buf0_), .Y(_4390_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_4330_), .B(_4390_), .Y(_4391_) );
INVX2 INVX2_151 ( .gnd(gnd), .vdd(vdd), .A(_4391_), .Y(module_0_W_182_) );
XNOR2X1 XNOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .B(bloque_datos_79_bF_buf1_), .Y(_4392_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_4332_), .B(_4392_), .Y(_4393_) );
INVX2 INVX2_152 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .Y(module_0_W_183_) );
XNOR2X1 XNOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf0_), .B(bloque_datos_40_bF_buf4_), .Y(_4394_) );
NAND3X1 NAND3X1_965 ( .gnd(gnd), .vdd(vdd), .A(_4335_), .B(_4394_), .C(_4334_), .Y(module_0_W_184_) );
XNOR2X1 XNOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf0_), .B(bloque_datos_41_bF_buf3_), .Y(_4395_) );
NAND3X1 NAND3X1_966 ( .gnd(gnd), .vdd(vdd), .A(_4340_), .B(_4395_), .C(_4339_), .Y(module_0_W_185_) );
XNOR2X1 XNOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf0_), .B(bloque_datos_42_bF_buf3_), .Y(_4396_) );
NAND3X1 NAND3X1_967 ( .gnd(gnd), .vdd(vdd), .A(_4343_), .B(_4396_), .C(_4342_), .Y(module_0_W_186_) );
XNOR2X1 XNOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf0_), .B(bloque_datos_43_bF_buf3_), .Y(_4397_) );
NAND3X1 NAND3X1_968 ( .gnd(gnd), .vdd(vdd), .A(_4346_), .B(_4397_), .C(_4345_), .Y(module_0_W_187_) );
XNOR2X1 XNOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf0_), .B(bloque_datos_44_bF_buf4_), .Y(_4398_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_4348_), .B(_4398_), .Y(_4399_) );
INVX1 INVX1_624 ( .gnd(gnd), .vdd(vdd), .A(_4399_), .Y(module_0_W_188_) );
XNOR2X1 XNOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf0_), .B(bloque_datos_45_bF_buf4_), .Y(_4400_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_4350_), .B(_4400_), .Y(_4401_) );
INVX1 INVX1_625 ( .gnd(gnd), .vdd(vdd), .A(_4401_), .Y(module_0_W_189_) );
XNOR2X1 XNOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf0_), .B(bloque_datos_46_bF_buf4_), .Y(_4402_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_4352_), .B(_4402_), .Y(_4403_) );
INVX1 INVX1_626 ( .gnd(gnd), .vdd(vdd), .A(_4403_), .Y(module_0_W_190_) );
XNOR2X1 XNOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf0_), .B(bloque_datos_47_bF_buf0_), .Y(_4404_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_4354_), .B(_4404_), .Y(_4405_) );
INVX1 INVX1_627 ( .gnd(gnd), .vdd(vdd), .A(_4405_), .Y(module_0_W_191_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf0_), .B(bloque_datos_48_bF_buf0_), .Y(_4406_) );
NOR2X1 NOR2X1_344 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf4_), .B(bloque_datos_48_bF_buf4_), .Y(_4407_) );
OAI21X1 OAI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_4406_), .B(_4407_), .C(_4356_), .Y(module_0_W_192_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf1_), .B(bloque_datos_49_bF_buf1_), .Y(_4408_) );
NOR2X1 NOR2X1_345 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf0_), .B(bloque_datos_49_bF_buf0_), .Y(_4409_) );
OAI21X1 OAI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(_4408_), .B(_4409_), .C(_4358_), .Y(module_0_W_193_) );
AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf0_), .B(bloque_datos_50_bF_buf0_), .Y(_4410_) );
NOR2X1 NOR2X1_346 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf4_), .B(bloque_datos_50_bF_buf3_), .Y(_4411_) );
OAI21X1 OAI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_4410_), .B(_4411_), .C(_4360_), .Y(module_0_W_194_) );
OR2X2 OR2X2_90 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_171_), .B(bloque_datos_51_bF_buf4_), .Y(module_0_W_195_) );
NOR2X1 NOR2X1_347 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf4_), .B(module_0_W_172_), .Y(_4412_) );
INVX1 INVX1_628 ( .gnd(gnd), .vdd(vdd), .A(_4412_), .Y(module_0_W_196_) );
NOR2X1 NOR2X1_348 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf3_), .B(module_0_W_173_), .Y(_4413_) );
INVX1 INVX1_629 ( .gnd(gnd), .vdd(vdd), .A(_4413_), .Y(module_0_W_197_) );
OR2X2 OR2X2_91 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_174_), .B(bloque_datos_54_bF_buf3_), .Y(module_0_W_198_) );
XNOR2X1 XNOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf0_), .B(bloque_datos[55]), .Y(_4414_) );
NAND2X1 NAND2X1_628 ( .gnd(gnd), .vdd(vdd), .A(_4414_), .B(_4373_), .Y(module_0_W_199_) );
NAND2X1 NAND2X1_629 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf0_), .B(module_0_W_128_), .Y(_4415_) );
INVX1 INVX1_630 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf4_), .Y(_4416_) );
NAND2X1 NAND2X1_630 ( .gnd(gnd), .vdd(vdd), .A(_4416_), .B(_4313_), .Y(_4417_) );
AOI21X1 AOI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_4417_), .B(_4415_), .C(module_0_W_176_), .Y(_4418_) );
INVX2 INVX2_153 ( .gnd(gnd), .vdd(vdd), .A(_4418_), .Y(module_0_W_200_) );
NAND2X1 NAND2X1_631 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf0_), .B(module_0_W_129_), .Y(_4419_) );
OR2X2 OR2X2_92 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_129_), .B(bloque_datos_57_bF_buf3_), .Y(_4420_) );
AOI21X1 AOI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_4419_), .B(_4420_), .C(module_0_W_177_), .Y(_4421_) );
INVX1 INVX1_631 ( .gnd(gnd), .vdd(vdd), .A(_4421_), .Y(module_0_W_201_) );
NAND2X1 NAND2X1_632 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf0_), .B(module_0_W_130_), .Y(_4422_) );
INVX1 INVX1_632 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf4_), .Y(_4423_) );
NAND2X1 NAND2X1_633 ( .gnd(gnd), .vdd(vdd), .A(_4423_), .B(_4317_), .Y(_4424_) );
AOI21X1 AOI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_4424_), .B(_4422_), .C(module_0_W_178_), .Y(_4425_) );
INVX1 INVX1_633 ( .gnd(gnd), .vdd(vdd), .A(_4425_), .Y(module_0_W_202_) );
NAND2X1 NAND2X1_634 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf0_), .B(module_0_W_131_), .Y(_4426_) );
INVX1 INVX1_634 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf4_), .Y(_4427_) );
NAND2X1 NAND2X1_635 ( .gnd(gnd), .vdd(vdd), .A(_4427_), .B(_4319_), .Y(_4428_) );
AOI21X1 AOI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_4428_), .B(_4426_), .C(module_0_W_179_), .Y(_4429_) );
INVX1 INVX1_635 ( .gnd(gnd), .vdd(vdd), .A(_4429_), .Y(module_0_W_203_) );
XNOR2X1 XNOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_132_), .B(bloque_datos_60_bF_buf3_), .Y(_4430_) );
NAND2X1 NAND2X1_636 ( .gnd(gnd), .vdd(vdd), .A(_4430_), .B(_4383_), .Y(module_0_W_204_) );
NAND2X1 NAND2X1_637 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf0_), .B(module_0_W_133_), .Y(_4431_) );
OR2X2 OR2X2_93 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_133_), .B(bloque_datos_61_bF_buf4_), .Y(_4432_) );
AOI21X1 AOI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_4431_), .B(_4432_), .C(module_0_W_181_), .Y(_4433_) );
INVX1 INVX1_636 ( .gnd(gnd), .vdd(vdd), .A(_4433_), .Y(module_0_W_205_) );
INVX2 INVX2_154 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf3_), .Y(_4434_) );
NAND2X1 NAND2X1_638 ( .gnd(gnd), .vdd(vdd), .A(_4434_), .B(_4391_), .Y(module_0_W_206_) );
INVX2 INVX2_155 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[63]), .Y(_4435_) );
NAND2X1 NAND2X1_639 ( .gnd(gnd), .vdd(vdd), .A(_4435_), .B(_4393_), .Y(module_0_W_207_) );
OAI21X1 OAI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(_4333_), .B(bloque_datos_80_bF_buf5_), .C(bloque_datos_64_bF_buf0_), .Y(_4436_) );
OR2X2 OR2X2_94 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_136_), .B(bloque_datos_64_bF_buf4_), .Y(_4437_) );
AOI21X1 AOI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_4436_), .B(_4437_), .C(module_0_W_184_), .Y(_4438_) );
INVX1 INVX1_637 ( .gnd(gnd), .vdd(vdd), .A(_4438_), .Y(module_0_W_208_) );
NAND2X1 NAND2X1_640 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_65_bF_buf0_), .B(module_0_W_137_), .Y(_4439_) );
OR2X2 OR2X2_95 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_137_), .B(bloque_datos_65_bF_buf3_), .Y(_4440_) );
AOI21X1 AOI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_4439_), .B(_4440_), .C(module_0_W_185_), .Y(_4441_) );
INVX1 INVX1_638 ( .gnd(gnd), .vdd(vdd), .A(_4441_), .Y(module_0_W_209_) );
OAI21X1 OAI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_4341_), .B(bloque_datos_82_bF_buf4_), .C(bloque_datos_66_bF_buf0_), .Y(_4442_) );
OR2X2 OR2X2_96 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_138_), .B(bloque_datos_66_bF_buf4_), .Y(_4443_) );
AOI21X1 AOI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_4442_), .B(_4443_), .C(module_0_W_186_), .Y(_4444_) );
INVX1 INVX1_639 ( .gnd(gnd), .vdd(vdd), .A(_4444_), .Y(module_0_W_210_) );
OAI21X1 OAI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(_4344_), .B(bloque_datos_83_bF_buf5_), .C(bloque_datos_67_bF_buf4_), .Y(_4445_) );
OR2X2 OR2X2_97 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_139_), .B(bloque_datos_67_bF_buf3_), .Y(_4446_) );
AOI21X1 AOI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_4445_), .B(_4446_), .C(module_0_W_187_), .Y(_4447_) );
INVX1 INVX1_640 ( .gnd(gnd), .vdd(vdd), .A(_4447_), .Y(module_0_W_211_) );
NAND2X1 NAND2X1_641 ( .gnd(gnd), .vdd(vdd), .A(_4363_), .B(_4399_), .Y(module_0_W_212_) );
NAND2X1 NAND2X1_642 ( .gnd(gnd), .vdd(vdd), .A(_4366_), .B(_4401_), .Y(module_0_W_213_) );
NAND2X1 NAND2X1_643 ( .gnd(gnd), .vdd(vdd), .A(_4369_), .B(_4403_), .Y(module_0_W_214_) );
INVX1 INVX1_641 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf0_), .Y(_4448_) );
NAND2X1 NAND2X1_644 ( .gnd(gnd), .vdd(vdd), .A(_4448_), .B(_4405_), .Y(module_0_W_215_) );
OR2X2 OR2X2_98 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_192_), .B(bloque_datos_72_bF_buf4_), .Y(module_0_W_216_) );
OR2X2 OR2X2_99 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_193_), .B(bloque_datos_73_bF_buf0_), .Y(module_0_W_217_) );
OR2X2 OR2X2_100 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_194_), .B(bloque_datos_74_bF_buf4_), .Y(module_0_W_218_) );
OR2X2 OR2X2_101 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_195_), .B(bloque_datos_75_bF_buf3_), .Y(module_0_W_219_) );
NAND2X1 NAND2X1_645 ( .gnd(gnd), .vdd(vdd), .A(_4322_), .B(_4412_), .Y(module_0_W_220_) );
NAND2X1 NAND2X1_646 ( .gnd(gnd), .vdd(vdd), .A(_4385_), .B(_4413_), .Y(module_0_W_221_) );
OR2X2 OR2X2_102 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_198_), .B(bloque_datos_78_bF_buf4_), .Y(module_0_W_222_) );
OR2X2 OR2X2_103 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_199_), .B(bloque_datos_79_bF_buf0_), .Y(module_0_W_223_) );
XNOR2X1 XNOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_152_), .B(bloque_datos_80_bF_buf4_), .Y(_4449_) );
NAND2X1 NAND2X1_647 ( .gnd(gnd), .vdd(vdd), .A(_4418_), .B(_4449_), .Y(module_0_W_224_) );
OAI21X1 OAI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_129_), .B(_4315_), .C(bloque_datos_81_bF_buf4_), .Y(_4450_) );
NAND3X1 NAND3X1_969 ( .gnd(gnd), .vdd(vdd), .A(_4337_), .B(_4378_), .C(_4377_), .Y(_4451_) );
NAND2X1 NAND2X1_648 ( .gnd(gnd), .vdd(vdd), .A(_4450_), .B(_4451_), .Y(_4452_) );
NAND2X1 NAND2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_4452_), .B(_4421_), .Y(module_0_W_225_) );
XNOR2X1 XNOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_154_), .B(bloque_datos_82_bF_buf3_), .Y(_4453_) );
NAND2X1 NAND2X1_650 ( .gnd(gnd), .vdd(vdd), .A(_4425_), .B(_4453_), .Y(module_0_W_226_) );
XNOR2X1 XNOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_155_), .B(bloque_datos_83_bF_buf4_), .Y(_4454_) );
NAND2X1 NAND2X1_651 ( .gnd(gnd), .vdd(vdd), .A(_4429_), .B(_4454_), .Y(module_0_W_227_) );
INVX1 INVX1_642 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf4_), .Y(_4455_) );
NAND3X1 NAND3X1_970 ( .gnd(gnd), .vdd(vdd), .A(_4455_), .B(_4430_), .C(_4383_), .Y(module_0_W_228_) );
OAI21X1 OAI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_133_), .B(_4327_), .C(bloque_datos_85_bF_buf4_), .Y(_4456_) );
INVX1 INVX1_643 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf3_), .Y(_4457_) );
NAND3X1 NAND3X1_971 ( .gnd(gnd), .vdd(vdd), .A(_4457_), .B(_4388_), .C(_4387_), .Y(_4458_) );
NAND2X1 NAND2X1_652 ( .gnd(gnd), .vdd(vdd), .A(_4456_), .B(_4458_), .Y(_4459_) );
NAND2X1 NAND2X1_653 ( .gnd(gnd), .vdd(vdd), .A(_4459_), .B(_4433_), .Y(module_0_W_229_) );
INVX1 INVX1_644 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf4_), .Y(_4460_) );
NAND3X1 NAND3X1_972 ( .gnd(gnd), .vdd(vdd), .A(_4460_), .B(_4434_), .C(_4391_), .Y(module_0_W_230_) );
INVX1 INVX1_645 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf3_), .Y(_4461_) );
NAND3X1 NAND3X1_973 ( .gnd(gnd), .vdd(vdd), .A(_4461_), .B(_4435_), .C(_4393_), .Y(module_0_W_231_) );
AOI21X1 AOI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_4335_), .B(_4334_), .C(_4282_), .Y(_4462_) );
NOR2X1 NOR2X1_349 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf3_), .B(module_0_W_160_), .Y(_4463_) );
OAI21X1 OAI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_4463_), .B(_4462_), .C(_4438_), .Y(module_0_W_232_) );
AOI21X1 AOI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_4340_), .B(_4339_), .C(_4286_), .Y(_4464_) );
NOR2X1 NOR2X1_350 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf3_), .B(module_0_W_161_), .Y(_4465_) );
OAI21X1 OAI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(_4464_), .B(_4465_), .C(_4441_), .Y(module_0_W_233_) );
AOI21X1 AOI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_4343_), .B(_4342_), .C(_4290_), .Y(_4466_) );
NOR2X1 NOR2X1_351 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf3_), .B(module_0_W_162_), .Y(_4467_) );
OAI21X1 OAI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(_4467_), .B(_4466_), .C(_4444_), .Y(module_0_W_234_) );
AOI21X1 AOI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_4346_), .B(_4345_), .C(_4294_), .Y(_4468_) );
NOR2X1 NOR2X1_352 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf3_), .B(module_0_W_163_), .Y(_4469_) );
OAI21X1 OAI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_4469_), .B(_4468_), .C(_4447_), .Y(module_0_W_235_) );
NAND3X1 NAND3X1_974 ( .gnd(gnd), .vdd(vdd), .A(_4298_), .B(_4363_), .C(_4399_), .Y(module_0_W_236_) );
NAND3X1 NAND3X1_975 ( .gnd(gnd), .vdd(vdd), .A(_4302_), .B(_4366_), .C(_4401_), .Y(module_0_W_237_) );
NAND3X1 NAND3X1_976 ( .gnd(gnd), .vdd(vdd), .A(_4306_), .B(_4369_), .C(_4403_), .Y(module_0_W_238_) );
NAND3X1 NAND3X1_977 ( .gnd(gnd), .vdd(vdd), .A(_4310_), .B(_4448_), .C(_4405_), .Y(module_0_W_239_) );
OR2X2 OR2X2_104 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_192_), .B(module_0_W_128_), .Y(module_0_W_240_) );
OR2X2 OR2X2_105 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_193_), .B(module_0_W_129_), .Y(module_0_W_241_) );
OR2X2 OR2X2_106 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_194_), .B(module_0_W_130_), .Y(module_0_W_242_) );
OR2X2 OR2X2_107 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_195_), .B(module_0_W_131_), .Y(module_0_W_243_) );
NAND2X1 NAND2X1_654 ( .gnd(gnd), .vdd(vdd), .A(_4324_), .B(_4412_), .Y(module_0_W_244_) );
NAND2X1 NAND2X1_655 ( .gnd(gnd), .vdd(vdd), .A(_4387_), .B(_4413_), .Y(module_0_W_245_) );
OR2X2 OR2X2_108 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_198_), .B(module_0_W_134_), .Y(module_0_W_246_) );
OR2X2 OR2X2_109 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_199_), .B(module_0_W_135_), .Y(module_0_W_247_) );
XNOR2X1 XNOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_176_), .B(module_0_W_136_), .Y(_4470_) );
NAND3X1 NAND3X1_978 ( .gnd(gnd), .vdd(vdd), .A(_4418_), .B(_4449_), .C(_4470_), .Y(module_0_W_248_) );
NAND3X1 NAND3X1_979 ( .gnd(gnd), .vdd(vdd), .A(_4339_), .B(_4452_), .C(_4421_), .Y(module_0_W_249_) );
XNOR2X1 XNOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_178_), .B(module_0_W_138_), .Y(_4471_) );
NAND3X1 NAND3X1_980 ( .gnd(gnd), .vdd(vdd), .A(_4425_), .B(_4453_), .C(_4471_), .Y(module_0_W_250_) );
XNOR2X1 XNOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_179_), .B(module_0_W_139_), .Y(_4472_) );
NAND3X1 NAND3X1_981 ( .gnd(gnd), .vdd(vdd), .A(_4429_), .B(_4454_), .C(_4472_), .Y(module_0_W_251_) );
INVX1 INVX1_646 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_140_), .Y(_4473_) );
NAND3X1 NAND3X1_982 ( .gnd(gnd), .vdd(vdd), .A(_4473_), .B(_4430_), .C(_4383_), .Y(module_0_W_252_) );
INVX1 INVX1_647 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_141_), .Y(_4474_) );
NAND3X1 NAND3X1_983 ( .gnd(gnd), .vdd(vdd), .A(_4474_), .B(_4459_), .C(_4433_), .Y(module_0_W_253_) );
INVX1 INVX1_648 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_142_), .Y(_4475_) );
NAND3X1 NAND3X1_984 ( .gnd(gnd), .vdd(vdd), .A(_4434_), .B(_4475_), .C(_4391_), .Y(module_0_W_254_) );
INVX1 INVX1_649 ( .gnd(gnd), .vdd(vdd), .A(module_0_W_143_), .Y(_4476_) );
NAND3X1 NAND3X1_985 ( .gnd(gnd), .vdd(vdd), .A(_4435_), .B(_4476_), .C(_4393_), .Y(module_0_W_255_) );
NAND3X1 NAND3X1_986 ( .gnd(gnd), .vdd(vdd), .A(_4709_), .B(_4710_), .C(_4711_), .Y(_4712_) );
NAND2X1 NAND2X1_656 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_200_), .B(_4694_), .Y(_4713_) );
OR2X2 OR2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_4694_), .B(module_1_W_200_), .Y(_4714_) );
NAND2X1 NAND2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_4713_), .B(_4714_), .Y(_4715_) );
NAND3X1 NAND3X1_987 ( .gnd(gnd), .vdd(vdd), .A(_4712_), .B(_4715_), .C(_4707_), .Y(_4716_) );
NAND2X1 NAND2X1_658 ( .gnd(gnd), .vdd(vdd), .A(_4712_), .B(_4707_), .Y(_4717_) );
INVX2 INVX2_156 ( .gnd(gnd), .vdd(vdd), .A(_4715_), .Y(_4718_) );
AOI21X1 AOI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_4718_), .B(_4717_), .C(_6700_), .Y(_4719_) );
NAND3X1 NAND3X1_988 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_228_), .B(_4716_), .C(_4719_), .Y(_4720_) );
INVX1 INVX1_650 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_228_), .Y(_4721_) );
AOI21X1 AOI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_4710_), .B(_4711_), .C(_4709_), .Y(_4722_) );
NAND3X1 NAND3X1_989 ( .gnd(gnd), .vdd(vdd), .A(_8129_), .B(_4702_), .C(_4699_), .Y(_4723_) );
NAND3X1 NAND3X1_990 ( .gnd(gnd), .vdd(vdd), .A(_8132_), .B(_4704_), .C(_4705_), .Y(_4724_) );
AOI21X1 AOI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_4723_), .B(_4724_), .C(_8185_), .Y(_4725_) );
OAI21X1 OAI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(_4722_), .B(_4725_), .C(_4718_), .Y(_4726_) );
NAND3X1 NAND3X1_991 ( .gnd(gnd), .vdd(vdd), .A(_6689_), .B(_4716_), .C(_4726_), .Y(_4727_) );
NAND2X1 NAND2X1_659 ( .gnd(gnd), .vdd(vdd), .A(_4721_), .B(_4727_), .Y(_4728_) );
AOI21X1 AOI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_4728_), .B(_4720_), .C(_8141_), .Y(_4729_) );
INVX1 INVX1_651 ( .gnd(gnd), .vdd(vdd), .A(_8141_), .Y(_4730_) );
NAND2X1 NAND2X1_660 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_228_), .B(_4727_), .Y(_4731_) );
NAND3X1 NAND3X1_992 ( .gnd(gnd), .vdd(vdd), .A(_4721_), .B(_4716_), .C(_4719_), .Y(_4732_) );
AOI21X1 AOI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(_4731_), .B(_4732_), .C(_4730_), .Y(_4733_) );
OAI21X1 OAI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_4729_), .B(_4733_), .C(_8183_), .Y(_4734_) );
OAI21X1 OAI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(_8147_), .B(_8149_), .C(_8142_), .Y(_4735_) );
NAND3X1 NAND3X1_993 ( .gnd(gnd), .vdd(vdd), .A(_4730_), .B(_4731_), .C(_4732_), .Y(_4736_) );
NAND3X1 NAND3X1_994 ( .gnd(gnd), .vdd(vdd), .A(_8141_), .B(_4728_), .C(_4720_), .Y(_4737_) );
NAND3X1 NAND3X1_995 ( .gnd(gnd), .vdd(vdd), .A(_4735_), .B(_4736_), .C(_4737_), .Y(_4738_) );
NAND2X1 NAND2X1_661 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_216_), .B(_4715_), .Y(_4739_) );
OR2X2 OR2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_4715_), .B(module_1_W_216_), .Y(_4740_) );
NAND2X1 NAND2X1_662 ( .gnd(gnd), .vdd(vdd), .A(_4739_), .B(_4740_), .Y(_4741_) );
NAND3X1 NAND3X1_996 ( .gnd(gnd), .vdd(vdd), .A(_4738_), .B(_4741_), .C(_4734_), .Y(_4742_) );
AOI21X1 AOI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_4736_), .B(_4737_), .C(_4735_), .Y(_4743_) );
NOR3X1 NOR3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_4729_), .B(_4733_), .C(_8183_), .Y(_4744_) );
INVX2 INVX2_157 ( .gnd(gnd), .vdd(vdd), .A(_4741_), .Y(_4745_) );
OAI21X1 OAI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_4744_), .B(_4743_), .C(_4745_), .Y(_4746_) );
NAND3X1 NAND3X1_997 ( .gnd(gnd), .vdd(vdd), .A(_7934_), .B(_4742_), .C(_4746_), .Y(_4747_) );
NAND2X1 NAND2X1_663 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_244_), .B(_4747_), .Y(_4748_) );
INVX1 INVX1_652 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_244_), .Y(_4749_) );
NAND2X1 NAND2X1_664 ( .gnd(gnd), .vdd(vdd), .A(_4738_), .B(_4734_), .Y(_4750_) );
AOI21X1 AOI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_4745_), .B(_4750_), .C(_7935_), .Y(_4751_) );
NAND3X1 NAND3X1_998 ( .gnd(gnd), .vdd(vdd), .A(_4749_), .B(_4742_), .C(_4751_), .Y(_4752_) );
NAND3X1 NAND3X1_999 ( .gnd(gnd), .vdd(vdd), .A(_8182_), .B(_4752_), .C(_4748_), .Y(_4753_) );
NAND3X1 NAND3X1_1000 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_244_), .B(_4742_), .C(_4751_), .Y(_4754_) );
NAND2X1 NAND2X1_665 ( .gnd(gnd), .vdd(vdd), .A(_4749_), .B(_4747_), .Y(_4755_) );
NAND3X1 NAND3X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_8154_), .B(_4754_), .C(_4755_), .Y(_4756_) );
AOI21X1 AOI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_4753_), .B(_4756_), .C(_8181_), .Y(_4757_) );
NOR2X1 NOR2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_7930_), .B(_8155_), .Y(_4758_) );
AOI21X1 AOI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_7945_), .B(_8158_), .C(_4758_), .Y(_4759_) );
AOI21X1 AOI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_4754_), .B(_4755_), .C(_8154_), .Y(_4760_) );
AOI21X1 AOI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_4752_), .B(_4748_), .C(_8182_), .Y(_4761_) );
NOR3X1 NOR3X1_135 ( .gnd(gnd), .vdd(vdd), .A(_4760_), .B(_4759_), .C(_4761_), .Y(_4762_) );
NOR2X1 NOR2X1_354 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_232_), .B(_4745_), .Y(_4763_) );
AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_4745_), .B(module_1_W_232_), .Y(_4764_) );
NOR2X1 NOR2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_4763_), .B(_4764_), .Y(_4765_) );
OAI21X1 OAI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(_4762_), .B(_4757_), .C(_4765_), .Y(_4766_) );
OAI21X1 OAI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_4760_), .B(_4761_), .C(_4759_), .Y(_4767_) );
NAND3X1 NAND3X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_4753_), .B(_4756_), .C(_8181_), .Y(_4768_) );
INVX2 INVX2_158 ( .gnd(gnd), .vdd(vdd), .A(_4765_), .Y(_4769_) );
NAND3X1 NAND3X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_4769_), .B(_4768_), .C(_4767_), .Y(_4770_) );
NAND2X1 NAND2X1_666 ( .gnd(gnd), .vdd(vdd), .A(_4770_), .B(_4766_), .Y(_4771_) );
XNOR2X1 XNOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_4771_), .B(_8178_), .Y(module_1_H_4_) );
NAND3X1 NAND3X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_8178_), .B(_4770_), .C(_4766_), .Y(_4772_) );
NOR2X1 NOR2X1_356 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_216_), .B(_4718_), .Y(_4773_) );
NOR2X1 NOR2X1_357 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_200_), .B(_4695_), .Y(_4774_) );
NOR2X1 NOR2X1_358 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_184_), .B(_4670_), .Y(_4775_) );
INVX1 INVX1_653 ( .gnd(gnd), .vdd(vdd), .A(_4648_), .Y(_4776_) );
NOR2X1 NOR2X1_359 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_168_), .B(_4776_), .Y(_4777_) );
NOR2X1 NOR2X1_360 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_152_), .B(_4626_), .Y(_4778_) );
INVX1 INVX1_654 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_153_), .Y(_4779_) );
NOR2X1 NOR2X1_361 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_136_), .B(_4603_), .Y(_4780_) );
INVX1 INVX1_655 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_137_), .Y(_4781_) );
INVX1 INVX1_656 ( .gnd(gnd), .vdd(vdd), .A(_4573_), .Y(_4782_) );
NOR2X1 NOR2X1_362 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf2_), .B(_4782_), .Y(_4783_) );
INVX1 INVX1_657 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf2_), .Y(_4784_) );
INVX1 INVX1_658 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_73_bF_buf3_), .Y(_4785_) );
NOR2X1 NOR2X1_363 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf3_), .B(_4523_), .Y(_4786_) );
NOR2X1 NOR2X1_364 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf3_), .B(_4498_), .Y(_4787_) );
NOR2X1 NOR2X1_365 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf3_), .B(_8284_), .Y(_4788_) );
NOR2X1 NOR2X1_366 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .B(_8259_), .Y(_4789_) );
INVX1 INVX1_659 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_25_), .Y(_4790_) );
INVX2 INVX2_159 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_9_), .Y(_4791_) );
NOR2X1 NOR2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_4790_), .B(_4791_), .Y(_4792_) );
NOR2X1 NOR2X1_368 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_25_), .B(module_1_W_9_), .Y(_4793_) );
NOR2X1 NOR2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_4793_), .B(_4792_), .Y(_4794_) );
NOR2X1 NOR2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_8257_), .B(_4794_), .Y(_4795_) );
AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_4794_), .B(_8257_), .Y(_4796_) );
NOR2X1 NOR2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_4795_), .B(_4796_), .Y(_4797_) );
NOR2X1 NOR2X1_372 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .B(_4797_), .Y(_4798_) );
INVX1 INVX1_660 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .Y(_4799_) );
OR2X2 OR2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_4796_), .B(_4795_), .Y(_4800_) );
NOR2X1 NOR2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_4799_), .B(_4800_), .Y(_4801_) );
OAI21X1 OAI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(_4801_), .B(_4798_), .C(_4789_), .Y(_4802_) );
OR2X2 OR2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_4801_), .B(_4798_), .Y(_4803_) );
OR2X2 OR2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_4803_), .B(_4789_), .Y(_4804_) );
AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_4804_), .B(_4802_), .Y(_4805_) );
NOR2X1 NOR2X1_374 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf2_), .B(_4805_), .Y(_4806_) );
AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_4805_), .B(bloque_datos_25_bF_buf1_), .Y(_4807_) );
OAI21X1 OAI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(_4807_), .B(_4806_), .C(_4788_), .Y(_4808_) );
OR2X2 OR2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_4807_), .B(_4806_), .Y(_4809_) );
OR2X2 OR2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_4809_), .B(_4788_), .Y(_4810_) );
AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_4810_), .B(_4808_), .Y(_4811_) );
NOR2X1 NOR2X1_375 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf2_), .B(_4811_), .Y(_4812_) );
INVX1 INVX1_661 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf1_), .Y(_4813_) );
NAND2X1 NAND2X1_667 ( .gnd(gnd), .vdd(vdd), .A(_4808_), .B(_4810_), .Y(_4814_) );
NOR2X1 NOR2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_4813_), .B(_4814_), .Y(_4815_) );
OAI21X1 OAI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_4812_), .B(_4815_), .C(_4787_), .Y(_4816_) );
OR2X2 OR2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_4812_), .B(_4815_), .Y(_4817_) );
OR2X2 OR2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_4817_), .B(_4787_), .Y(_4818_) );
AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_4818_), .B(_4816_), .Y(_4819_) );
NOR2X1 NOR2X1_377 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf2_), .B(_4819_), .Y(_4820_) );
INVX1 INVX1_662 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf1_), .Y(_4821_) );
NAND2X1 NAND2X1_668 ( .gnd(gnd), .vdd(vdd), .A(_4816_), .B(_4818_), .Y(_4822_) );
NOR2X1 NOR2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_4821_), .B(_4822_), .Y(_4823_) );
OAI21X1 OAI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_4820_), .B(_4823_), .C(_4786_), .Y(_4824_) );
OR2X2 OR2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_4820_), .B(_4823_), .Y(_4825_) );
OR2X2 OR2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_4825_), .B(_4786_), .Y(_4826_) );
NAND2X1 NAND2X1_669 ( .gnd(gnd), .vdd(vdd), .A(_4824_), .B(_4826_), .Y(_4827_) );
NAND2X1 NAND2X1_670 ( .gnd(gnd), .vdd(vdd), .A(_4785_), .B(_4827_), .Y(_4828_) );
OR2X2 OR2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_4827_), .B(_4785_), .Y(_4829_) );
NAND2X1 NAND2X1_671 ( .gnd(gnd), .vdd(vdd), .A(_4828_), .B(_4829_), .Y(_4830_) );
NAND2X1 NAND2X1_672 ( .gnd(gnd), .vdd(vdd), .A(_4570_), .B(_4830_), .Y(_4831_) );
OR2X2 OR2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_4830_), .B(_4570_), .Y(_4832_) );
NAND2X1 NAND2X1_673 ( .gnd(gnd), .vdd(vdd), .A(_4831_), .B(_4832_), .Y(_4833_) );
NAND2X1 NAND2X1_674 ( .gnd(gnd), .vdd(vdd), .A(_4784_), .B(_4833_), .Y(_4834_) );
OR2X2 OR2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_4833_), .B(_4784_), .Y(_4835_) );
NAND2X1 NAND2X1_675 ( .gnd(gnd), .vdd(vdd), .A(_4834_), .B(_4835_), .Y(_4836_) );
NAND2X1 NAND2X1_676 ( .gnd(gnd), .vdd(vdd), .A(_4783_), .B(_4836_), .Y(_4837_) );
NOR2X1 NOR2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_4783_), .B(_4836_), .Y(_4838_) );
INVX1 INVX1_663 ( .gnd(gnd), .vdd(vdd), .A(_4838_), .Y(_4839_) );
NAND2X1 NAND2X1_677 ( .gnd(gnd), .vdd(vdd), .A(_4837_), .B(_4839_), .Y(_4840_) );
NAND2X1 NAND2X1_678 ( .gnd(gnd), .vdd(vdd), .A(_4781_), .B(_4840_), .Y(_4841_) );
INVX2 INVX2_160 ( .gnd(gnd), .vdd(vdd), .A(_4840_), .Y(_4842_) );
NAND2X1 NAND2X1_679 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_137_), .B(_4842_), .Y(_4843_) );
NAND2X1 NAND2X1_680 ( .gnd(gnd), .vdd(vdd), .A(_4841_), .B(_4843_), .Y(_4844_) );
NAND2X1 NAND2X1_681 ( .gnd(gnd), .vdd(vdd), .A(_4780_), .B(_4844_), .Y(_4845_) );
NOR2X1 NOR2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_4780_), .B(_4844_), .Y(_4846_) );
INVX1 INVX1_664 ( .gnd(gnd), .vdd(vdd), .A(_4846_), .Y(_4847_) );
NAND2X1 NAND2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_4845_), .B(_4847_), .Y(_4848_) );
NAND2X1 NAND2X1_683 ( .gnd(gnd), .vdd(vdd), .A(_4779_), .B(_4848_), .Y(_4849_) );
NOR2X1 NOR2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_4779_), .B(_4848_), .Y(_4850_) );
INVX1 INVX1_665 ( .gnd(gnd), .vdd(vdd), .A(_4850_), .Y(_4851_) );
NAND2X1 NAND2X1_684 ( .gnd(gnd), .vdd(vdd), .A(_4849_), .B(_4851_), .Y(_4852_) );
NAND2X1 NAND2X1_685 ( .gnd(gnd), .vdd(vdd), .A(_4778_), .B(_4852_), .Y(_4853_) );
NOR2X1 NOR2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_4778_), .B(_4852_), .Y(_4854_) );
INVX1 INVX1_666 ( .gnd(gnd), .vdd(vdd), .A(_4854_), .Y(_4855_) );
NAND2X1 NAND2X1_686 ( .gnd(gnd), .vdd(vdd), .A(_4853_), .B(_4855_), .Y(_4856_) );
INVX2 INVX2_161 ( .gnd(gnd), .vdd(vdd), .A(_4856_), .Y(_4857_) );
NOR2X1 NOR2X1_383 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_169_), .B(_4857_), .Y(_4858_) );
NAND2X1 NAND2X1_687 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_169_), .B(_4857_), .Y(_4859_) );
INVX2 INVX2_162 ( .gnd(gnd), .vdd(vdd), .A(_4859_), .Y(_4860_) );
OAI21X1 OAI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_4860_), .B(_4858_), .C(_4777_), .Y(_4861_) );
NOR2X1 NOR2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_4858_), .B(_4860_), .Y(_4862_) );
OAI21X1 OAI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_168_), .B(_4776_), .C(_4862_), .Y(_4863_) );
NAND2X1 NAND2X1_688 ( .gnd(gnd), .vdd(vdd), .A(_4861_), .B(_4863_), .Y(_4864_) );
INVX2 INVX2_163 ( .gnd(gnd), .vdd(vdd), .A(_4864_), .Y(_4865_) );
NOR2X1 NOR2X1_385 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_185_), .B(_4865_), .Y(_4866_) );
NAND2X1 NAND2X1_689 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_185_), .B(_4865_), .Y(_4867_) );
INVX2 INVX2_164 ( .gnd(gnd), .vdd(vdd), .A(_4867_), .Y(_4868_) );
OAI21X1 OAI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_4868_), .B(_4866_), .C(_4775_), .Y(_4869_) );
NOR2X1 NOR2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_4866_), .B(_4868_), .Y(_4870_) );
OAI21X1 OAI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_184_), .B(_4670_), .C(_4870_), .Y(_4871_) );
NAND2X1 NAND2X1_690 ( .gnd(gnd), .vdd(vdd), .A(_4869_), .B(_4871_), .Y(_4872_) );
INVX2 INVX2_165 ( .gnd(gnd), .vdd(vdd), .A(_4872_), .Y(_4873_) );
NOR2X1 NOR2X1_387 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_201_), .B(_4873_), .Y(_4874_) );
NAND2X1 NAND2X1_691 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_201_), .B(_4873_), .Y(_4875_) );
INVX2 INVX2_166 ( .gnd(gnd), .vdd(vdd), .A(_4875_), .Y(_4876_) );
OAI21X1 OAI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_4876_), .B(_4874_), .C(_4774_), .Y(_4877_) );
NOR2X1 NOR2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_4874_), .B(_4876_), .Y(_4878_) );
OAI21X1 OAI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_200_), .B(_4695_), .C(_4878_), .Y(_4879_) );
NAND2X1 NAND2X1_692 ( .gnd(gnd), .vdd(vdd), .A(_4877_), .B(_4879_), .Y(_4880_) );
INVX2 INVX2_167 ( .gnd(gnd), .vdd(vdd), .A(_4880_), .Y(_4881_) );
NOR2X1 NOR2X1_389 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_217_), .B(_4881_), .Y(_4882_) );
NAND2X1 NAND2X1_693 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_217_), .B(_4881_), .Y(_4883_) );
INVX2 INVX2_168 ( .gnd(gnd), .vdd(vdd), .A(_4883_), .Y(_4884_) );
OAI21X1 OAI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_4884_), .B(_4882_), .C(_4773_), .Y(_4885_) );
NOR2X1 NOR2X1_390 ( .gnd(gnd), .vdd(vdd), .A(_4882_), .B(_4884_), .Y(_4886_) );
OAI21X1 OAI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_216_), .B(_4718_), .C(_4886_), .Y(_4887_) );
NAND2X1 NAND2X1_694 ( .gnd(gnd), .vdd(vdd), .A(_4885_), .B(_4887_), .Y(_4888_) );
INVX2 INVX2_169 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .Y(_4889_) );
NOR2X1 NOR2X1_391 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_233_), .B(_4889_), .Y(_4890_) );
NAND2X1 NAND2X1_695 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_233_), .B(_4889_), .Y(_4891_) );
INVX2 INVX2_170 ( .gnd(gnd), .vdd(vdd), .A(_4891_), .Y(_4892_) );
OAI21X1 OAI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_4892_), .B(_4890_), .C(_4763_), .Y(_4893_) );
NOR2X1 NOR2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_4890_), .B(_4892_), .Y(_4894_) );
OAI21X1 OAI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_232_), .B(_4745_), .C(_4894_), .Y(_4895_) );
NAND2X1 NAND2X1_696 ( .gnd(gnd), .vdd(vdd), .A(_4893_), .B(_4895_), .Y(_4896_) );
OAI21X1 OAI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_4761_), .B(_4759_), .C(_4753_), .Y(_4897_) );
INVX1 INVX1_667 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_245_), .Y(_4898_) );
AOI21X1 AOI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_4735_), .B(_4737_), .C(_4729_), .Y(_4899_) );
INVX2 INVX2_171 ( .gnd(gnd), .vdd(vdd), .A(_4731_), .Y(_4900_) );
INVX1 INVX1_668 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_229_), .Y(_4901_) );
AOI21X1 AOI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(_4709_), .B(_4711_), .C(_4703_), .Y(_4902_) );
INVX2 INVX2_172 ( .gnd(gnd), .vdd(vdd), .A(_4704_), .Y(_4903_) );
INVX1 INVX1_669 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_213_), .Y(_4904_) );
AOI21X1 AOI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_4689_), .B(_4687_), .C(_4679_), .Y(_4905_) );
INVX2 INVX2_173 ( .gnd(gnd), .vdd(vdd), .A(_4683_), .Y(_4906_) );
INVX1 INVX1_670 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_197_), .Y(_4907_) );
AOI21X1 AOI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_4663_), .B(_4661_), .C(_4656_), .Y(_4908_) );
INVX2 INVX2_174 ( .gnd(gnd), .vdd(vdd), .A(_4657_), .Y(_4909_) );
INVX1 INVX1_671 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_181_), .Y(_4910_) );
AOI21X1 AOI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_8191_), .B(_4644_), .C(_4637_), .Y(_4911_) );
INVX2 INVX2_175 ( .gnd(gnd), .vdd(vdd), .A(_4639_), .Y(_4912_) );
INVX1 INVX1_672 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_165_), .Y(_4913_) );
INVX1 INVX1_673 ( .gnd(gnd), .vdd(vdd), .A(_4848_), .Y(_4914_) );
AOI21X1 AOI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(_4617_), .B(_4619_), .C(_4612_), .Y(_4915_) );
INVX1 INVX1_674 ( .gnd(gnd), .vdd(vdd), .A(_4613_), .Y(_4916_) );
INVX1 INVX1_675 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_149_), .Y(_4917_) );
AOI21X1 AOI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_4589_), .B(_8194_), .C(_4599_), .Y(_4918_) );
AOI21X1 AOI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(_4562_), .B(_4563_), .C(_8196_), .Y(_4919_) );
AOI21X1 AOI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_4566_), .B(_4568_), .C(_4919_), .Y(_4920_) );
NOR3X1 NOR3X1_136 ( .gnd(gnd), .vdd(vdd), .A(_4530_), .B(_8048_), .C(_4534_), .Y(_4921_) );
OAI21X1 OAI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_4921_), .B(_8198_), .C(_4543_), .Y(_4922_) );
AOI21X1 AOI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_4512_), .B(_4513_), .C(_8202_), .Y(_4923_) );
AOI21X1 AOI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_4518_), .B(_4516_), .C(_4923_), .Y(_4924_) );
AOI21X1 AOI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_4487_), .B(_4488_), .C(_8206_), .Y(_4925_) );
AOI21X1 AOI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_4493_), .B(_4491_), .C(_4925_), .Y(_4926_) );
INVX1 INVX1_676 ( .gnd(gnd), .vdd(vdd), .A(_8277_), .Y(_4927_) );
AOI21X1 AOI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_8276_), .B(_8278_), .C(_4927_), .Y(_4928_) );
INVX1 INVX1_677 ( .gnd(gnd), .vdd(vdd), .A(_8253_), .Y(_4929_) );
AOI21X1 AOI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_8254_), .B(_8252_), .C(_4929_), .Y(_4930_) );
AOI21X1 AOI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(_8226_), .B(_8225_), .C(_7985_), .Y(_4931_) );
NOR2X1 NOR2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .B(_8237_), .Y(_4932_) );
INVX1 INVX1_678 ( .gnd(gnd), .vdd(vdd), .A(_8225_), .Y(_4933_) );
NOR2X1 NOR2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_7084_), .B(_7073_), .Y(_4934_) );
INVX2 INVX2_176 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_5_), .Y(_4935_) );
XNOR2X1 XNOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_8217_), .B(_4935_), .Y(_4936_) );
NAND2X1 NAND2X1_697 ( .gnd(gnd), .vdd(vdd), .A(_4934_), .B(_4936_), .Y(_4937_) );
INVX1 INVX1_679 ( .gnd(gnd), .vdd(vdd), .A(_4934_), .Y(_4938_) );
NOR2X1 NOR2X1_395 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_5_), .B(_8217_), .Y(_4939_) );
NOR2X1 NOR2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_4935_), .B(_8214_), .Y(_4940_) );
OAI21X1 OAI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(_4940_), .B(_4939_), .C(_4938_), .Y(_4941_) );
NAND3X1 NAND3X1_1005 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_21_), .B(_4937_), .C(_4941_), .Y(_4942_) );
INVX1 INVX1_680 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_21_), .Y(_4943_) );
OAI21X1 OAI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_4940_), .B(_4939_), .C(_4934_), .Y(_4944_) );
OAI21X1 OAI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_7073_), .B(_7084_), .C(_4936_), .Y(_4945_) );
NAND3X1 NAND3X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_4943_), .B(_4945_), .C(_4944_), .Y(_4946_) );
NAND3X1 NAND3X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_4933_), .B(_4942_), .C(_4946_), .Y(_4947_) );
NAND3X1 NAND3X1_1008 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_21_), .B(_4945_), .C(_4944_), .Y(_4948_) );
NAND3X1 NAND3X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_4943_), .B(_4937_), .C(_4941_), .Y(_4949_) );
NAND3X1 NAND3X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_8225_), .B(_4949_), .C(_4948_), .Y(_4950_) );
AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_4947_), .B(_4950_), .Y(_4951_) );
NAND2X1 NAND2X1_698 ( .gnd(gnd), .vdd(vdd), .A(_4951_), .B(_4932_), .Y(_4952_) );
NAND2X1 NAND2X1_699 ( .gnd(gnd), .vdd(vdd), .A(_4950_), .B(_4947_), .Y(_4953_) );
OAI21X1 OAI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .B(_8237_), .C(_4953_), .Y(_4954_) );
XNOR2X1 XNOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_7160_), .B(module_1_W_9_), .Y(_4955_) );
NAND3X1 NAND3X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_4955_), .B(_4954_), .C(_4952_), .Y(_4956_) );
NAND2X1 NAND2X1_700 ( .gnd(gnd), .vdd(vdd), .A(_8224_), .B(_8228_), .Y(_4957_) );
NOR2X1 NOR2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_4953_), .B(_4957_), .Y(_4958_) );
NOR2X1 NOR2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_4951_), .B(_4932_), .Y(_4959_) );
INVX1 INVX1_681 ( .gnd(gnd), .vdd(vdd), .A(_4955_), .Y(_4960_) );
OAI21X1 OAI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_4959_), .B(_4958_), .C(_4960_), .Y(_4961_) );
NAND3X1 NAND3X1_1012 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf3_), .B(_4956_), .C(_4961_), .Y(_4962_) );
INVX1 INVX1_682 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf2_), .Y(_4963_) );
NAND3X1 NAND3X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_4960_), .B(_4954_), .C(_4952_), .Y(_4964_) );
OAI21X1 OAI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_4959_), .B(_4958_), .C(_4955_), .Y(_4965_) );
NAND3X1 NAND3X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_4963_), .B(_4964_), .C(_4965_), .Y(_4966_) );
NAND3X1 NAND3X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_8240_), .B(_4962_), .C(_4966_), .Y(_4967_) );
NAND3X1 NAND3X1_1016 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf1_), .B(_4964_), .C(_4965_), .Y(_4968_) );
NAND3X1 NAND3X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_4963_), .B(_4956_), .C(_4961_), .Y(_4969_) );
NAND3X1 NAND3X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_8246_), .B(_4968_), .C(_4969_), .Y(_4970_) );
NAND3X1 NAND3X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_4930_), .B(_4967_), .C(_4970_), .Y(_4971_) );
NAND2X1 NAND2X1_701 ( .gnd(gnd), .vdd(vdd), .A(_8253_), .B(_8255_), .Y(_4972_) );
NAND3X1 NAND3X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_8246_), .B(_4962_), .C(_4966_), .Y(_4973_) );
NAND3X1 NAND3X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_8240_), .B(_4968_), .C(_4969_), .Y(_4974_) );
NAND3X1 NAND3X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_4973_), .B(_4974_), .C(_4972_), .Y(_4975_) );
XNOR2X1 XNOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_7204_), .B(_4797_), .Y(_4976_) );
INVX1 INVX1_683 ( .gnd(gnd), .vdd(vdd), .A(_4976_), .Y(_4977_) );
NAND3X1 NAND3X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_4971_), .B(_4977_), .C(_4975_), .Y(_4978_) );
AOI21X1 AOI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_4973_), .B(_4974_), .C(_4972_), .Y(_4979_) );
AOI21X1 AOI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_4967_), .B(_4970_), .C(_4930_), .Y(_4980_) );
OAI21X1 OAI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_4979_), .B(_4980_), .C(_4976_), .Y(_4981_) );
NAND3X1 NAND3X1_1024 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf3_), .B(_4978_), .C(_4981_), .Y(_4982_) );
INVX1 INVX1_684 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf2_), .Y(_4983_) );
NAND3X1 NAND3X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_4971_), .B(_4976_), .C(_4975_), .Y(_4984_) );
OAI21X1 OAI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_4979_), .B(_4980_), .C(_4977_), .Y(_4985_) );
NAND3X1 NAND3X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_4983_), .B(_4984_), .C(_4985_), .Y(_4986_) );
NAND3X1 NAND3X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_8266_), .B(_4982_), .C(_4986_), .Y(_4987_) );
NAND3X1 NAND3X1_1028 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf1_), .B(_4984_), .C(_4985_), .Y(_4988_) );
NAND3X1 NAND3X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_4983_), .B(_4978_), .C(_4981_), .Y(_4989_) );
NAND3X1 NAND3X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_8272_), .B(_4988_), .C(_4989_), .Y(_4990_) );
NAND3X1 NAND3X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_4987_), .B(_4990_), .C(_4928_), .Y(_4991_) );
INVX1 INVX1_685 ( .gnd(gnd), .vdd(vdd), .A(_8278_), .Y(_4992_) );
OAI21X1 OAI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_4992_), .B(_8207_), .C(_8277_), .Y(_4993_) );
NAND3X1 NAND3X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_8272_), .B(_4982_), .C(_4986_), .Y(_4994_) );
NAND3X1 NAND3X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_8266_), .B(_4988_), .C(_4989_), .Y(_4995_) );
NAND3X1 NAND3X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_4994_), .B(_4993_), .C(_4995_), .Y(_4996_) );
NAND2X1 NAND2X1_702 ( .gnd(gnd), .vdd(vdd), .A(_4802_), .B(_4804_), .Y(_4997_) );
XNOR2X1 XNOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_7259_), .B(_4997_), .Y(_4998_) );
INVX1 INVX1_686 ( .gnd(gnd), .vdd(vdd), .A(_4998_), .Y(_4999_) );
NAND3X1 NAND3X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_4999_), .B(_4996_), .C(_4991_), .Y(_5000_) );
AOI21X1 AOI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_4994_), .B(_4995_), .C(_4993_), .Y(_5001_) );
AOI21X1 AOI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_4987_), .B(_4990_), .C(_4928_), .Y(_5002_) );
OAI21X1 OAI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_5001_), .B(_5002_), .C(_4998_), .Y(_5003_) );
NAND3X1 NAND3X1_1036 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf2_), .B(_5000_), .C(_5003_), .Y(_5004_) );
INVX1 INVX1_687 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf1_), .Y(_5005_) );
NAND3X1 NAND3X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_4998_), .B(_4996_), .C(_4991_), .Y(_5006_) );
OAI21X1 OAI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(_5001_), .B(_5002_), .C(_4999_), .Y(_5007_) );
NAND3X1 NAND3X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_5005_), .B(_5006_), .C(_5007_), .Y(_5008_) );
NAND3X1 NAND3X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_4481_), .B(_5004_), .C(_5008_), .Y(_5009_) );
NAND3X1 NAND3X1_1040 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf0_), .B(_5006_), .C(_5007_), .Y(_5010_) );
NAND3X1 NAND3X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_5005_), .B(_5000_), .C(_5003_), .Y(_5011_) );
NAND3X1 NAND3X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_4487_), .B(_5010_), .C(_5011_), .Y(_5012_) );
NAND3X1 NAND3X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_4926_), .B(_5009_), .C(_5012_), .Y(_5013_) );
NOR3X1 NOR3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_4481_), .B(_8024_), .C(_4485_), .Y(_5014_) );
OAI21X1 OAI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(_5014_), .B(_8205_), .C(_4492_), .Y(_5015_) );
NAND3X1 NAND3X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_4487_), .B(_5004_), .C(_5008_), .Y(_5016_) );
NAND3X1 NAND3X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_4481_), .B(_5010_), .C(_5011_), .Y(_5017_) );
NAND3X1 NAND3X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_5015_), .B(_5016_), .C(_5017_), .Y(_5018_) );
XNOR2X1 XNOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_4811_), .Y(_5019_) );
NAND3X1 NAND3X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_5019_), .B(_5013_), .C(_5018_), .Y(_5020_) );
AOI21X1 AOI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_5016_), .B(_5017_), .C(_5015_), .Y(_5021_) );
AOI21X1 AOI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_5009_), .B(_5012_), .C(_4926_), .Y(_5022_) );
INVX1 INVX1_688 ( .gnd(gnd), .vdd(vdd), .A(_5019_), .Y(_5023_) );
OAI21X1 OAI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_5021_), .B(_5022_), .C(_5023_), .Y(_5024_) );
NAND3X1 NAND3X1_1048 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf2_), .B(_5020_), .C(_5024_), .Y(_5025_) );
INVX1 INVX1_689 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf1_), .Y(_5026_) );
NAND3X1 NAND3X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_5023_), .B(_5013_), .C(_5018_), .Y(_5027_) );
OAI21X1 OAI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_5021_), .B(_5022_), .C(_5019_), .Y(_5028_) );
NAND3X1 NAND3X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_5026_), .B(_5027_), .C(_5028_), .Y(_5029_) );
NAND3X1 NAND3X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_4505_), .B(_5025_), .C(_5029_), .Y(_5030_) );
NAND3X1 NAND3X1_1052 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf0_), .B(_5027_), .C(_5028_), .Y(_5031_) );
NAND3X1 NAND3X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_5026_), .B(_5020_), .C(_5024_), .Y(_5032_) );
NAND3X1 NAND3X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_4512_), .B(_5031_), .C(_5032_), .Y(_5033_) );
NAND3X1 NAND3X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_4924_), .B(_5030_), .C(_5033_), .Y(_5034_) );
NOR3X1 NOR3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_4505_), .B(_4511_), .C(_4509_), .Y(_5035_) );
OAI21X1 OAI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(_5035_), .B(_8200_), .C(_4517_), .Y(_5036_) );
NAND3X1 NAND3X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_4512_), .B(_5025_), .C(_5029_), .Y(_5037_) );
NAND3X1 NAND3X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_4505_), .B(_5031_), .C(_5032_), .Y(_5038_) );
NAND3X1 NAND3X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_5037_), .B(_5038_), .C(_5036_), .Y(_5039_) );
XNOR2X1 XNOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_7402_), .B(_4819_), .Y(_5040_) );
INVX1 INVX1_690 ( .gnd(gnd), .vdd(vdd), .A(_5040_), .Y(_5041_) );
NAND3X1 NAND3X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_5041_), .B(_5034_), .C(_5039_), .Y(_5042_) );
AOI21X1 AOI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_5037_), .B(_5038_), .C(_5036_), .Y(_5043_) );
AOI21X1 AOI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_5030_), .B(_5033_), .C(_4924_), .Y(_5044_) );
OAI21X1 OAI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_5043_), .B(_5044_), .C(_5040_), .Y(_5045_) );
NAND3X1 NAND3X1_1060 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf2_), .B(_5042_), .C(_5045_), .Y(_5046_) );
INVX1 INVX1_691 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf1_), .Y(_5047_) );
NAND3X1 NAND3X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_5040_), .B(_5034_), .C(_5039_), .Y(_5048_) );
OAI21X1 OAI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_5043_), .B(_5044_), .C(_5041_), .Y(_5049_) );
NAND3X1 NAND3X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_5047_), .B(_5048_), .C(_5049_), .Y(_5050_) );
NAND3X1 NAND3X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_4536_), .B(_5046_), .C(_5050_), .Y(_5051_) );
NAND3X1 NAND3X1_1064 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf0_), .B(_5048_), .C(_5049_), .Y(_5052_) );
NAND3X1 NAND3X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_5047_), .B(_5042_), .C(_5045_), .Y(_5053_) );
NAND3X1 NAND3X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_4530_), .B(_5052_), .C(_5053_), .Y(_5054_) );
AOI21X1 AOI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_5051_), .B(_5054_), .C(_4922_), .Y(_5055_) );
AOI21X1 AOI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_4536_), .B(_4537_), .C(_8199_), .Y(_5056_) );
AOI21X1 AOI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_4542_), .B(_4544_), .C(_5056_), .Y(_5057_) );
NAND3X1 NAND3X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_4530_), .B(_5046_), .C(_5050_), .Y(_5058_) );
NAND3X1 NAND3X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_4536_), .B(_5052_), .C(_5053_), .Y(_5059_) );
AOI21X1 AOI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_5058_), .B(_5059_), .C(_5057_), .Y(_5060_) );
XNOR2X1 XNOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_7446_), .B(_4827_), .Y(_5061_) );
NOR3X1 NOR3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_5060_), .B(_5061_), .C(_5055_), .Y(_5062_) );
NAND3X1 NAND3X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_5057_), .B(_5058_), .C(_5059_), .Y(_5063_) );
NAND3X1 NAND3X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_5051_), .B(_5054_), .C(_4922_), .Y(_5064_) );
INVX1 INVX1_692 ( .gnd(gnd), .vdd(vdd), .A(_5061_), .Y(_5065_) );
AOI21X1 AOI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_5063_), .B(_5064_), .C(_5065_), .Y(_5066_) );
OAI21X1 OAI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(_5062_), .B(_5066_), .C(bloque_datos_85_bF_buf2_), .Y(_5067_) );
INVX1 INVX1_693 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf1_), .Y(_5068_) );
NAND3X1 NAND3X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_5065_), .B(_5063_), .C(_5064_), .Y(_5069_) );
OAI21X1 OAI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_5055_), .B(_5060_), .C(_5061_), .Y(_5070_) );
NAND3X1 NAND3X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_5068_), .B(_5069_), .C(_5070_), .Y(_5071_) );
NAND3X1 NAND3X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_4556_), .B(_5071_), .C(_5067_), .Y(_5072_) );
NAND3X1 NAND3X1_1074 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf0_), .B(_5069_), .C(_5070_), .Y(_5073_) );
OAI21X1 OAI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(_5062_), .B(_5066_), .C(_5068_), .Y(_5074_) );
NAND3X1 NAND3X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_4562_), .B(_5073_), .C(_5074_), .Y(_5075_) );
NAND3X1 NAND3X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_4920_), .B(_5072_), .C(_5075_), .Y(_5076_) );
NOR3X1 NOR3X1_140 ( .gnd(gnd), .vdd(vdd), .A(_4556_), .B(_8060_), .C(_4560_), .Y(_5077_) );
OAI21X1 OAI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_5077_), .B(_8195_), .C(_4567_), .Y(_5078_) );
NAND3X1 NAND3X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_4562_), .B(_5071_), .C(_5067_), .Y(_5079_) );
NAND3X1 NAND3X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_4556_), .B(_5073_), .C(_5074_), .Y(_5080_) );
NAND3X1 NAND3X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_5079_), .B(_5080_), .C(_5078_), .Y(_5081_) );
XNOR2X1 XNOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_7544_), .B(_4833_), .Y(_5082_) );
NAND3X1 NAND3X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_5076_), .C(_5081_), .Y(_5083_) );
AOI21X1 AOI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_5079_), .B(_5080_), .C(_5078_), .Y(_5084_) );
AOI21X1 AOI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(_5072_), .B(_5075_), .C(_4920_), .Y(_5085_) );
INVX1 INVX1_694 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .Y(_5086_) );
OAI21X1 OAI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(_5084_), .B(_5085_), .C(_5086_), .Y(_5087_) );
NAND3X1 NAND3X1_1081 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_133_), .B(_5083_), .C(_5087_), .Y(_5088_) );
INVX1 INVX1_695 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_133_), .Y(_5089_) );
NAND3X1 NAND3X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_5086_), .B(_5076_), .C(_5081_), .Y(_5090_) );
OAI21X1 OAI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(_5084_), .B(_5085_), .C(_5082_), .Y(_5091_) );
NAND3X1 NAND3X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_5089_), .B(_5090_), .C(_5091_), .Y(_5092_) );
AOI21X1 AOI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_5088_), .B(_5092_), .C(_4580_), .Y(_5093_) );
NAND3X1 NAND3X1_1084 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_133_), .B(_5090_), .C(_5091_), .Y(_5094_) );
NAND3X1 NAND3X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_5089_), .B(_5083_), .C(_5087_), .Y(_5095_) );
AOI21X1 AOI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_5095_), .C(_4587_), .Y(_5096_) );
OAI21X1 OAI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(_5093_), .B(_5096_), .C(_4918_), .Y(_5097_) );
OAI21X1 OAI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_4600_), .B(_4591_), .C(_4585_), .Y(_5098_) );
AOI21X1 AOI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_5088_), .B(_5092_), .C(_4587_), .Y(_5099_) );
AOI21X1 AOI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_5095_), .C(_4580_), .Y(_5100_) );
OAI21X1 OAI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_5099_), .B(_5100_), .C(_5098_), .Y(_5101_) );
NAND3X1 NAND3X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_4842_), .B(_5097_), .C(_5101_), .Y(_5102_) );
NAND3X1 NAND3X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_4587_), .B(_5094_), .C(_5095_), .Y(_5103_) );
NAND3X1 NAND3X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_4580_), .B(_5088_), .C(_5092_), .Y(_5104_) );
AOI21X1 AOI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_5103_), .B(_5104_), .C(_5098_), .Y(_5105_) );
NAND3X1 NAND3X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_4580_), .B(_5094_), .C(_5095_), .Y(_5106_) );
NAND3X1 NAND3X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_4587_), .B(_5088_), .C(_5092_), .Y(_5107_) );
AOI21X1 AOI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(_5107_), .C(_4918_), .Y(_5108_) );
OAI21X1 OAI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .B(_5108_), .C(_4840_), .Y(_5109_) );
NAND2X1 NAND2X1_703 ( .gnd(gnd), .vdd(vdd), .A(_5102_), .B(_5109_), .Y(_5110_) );
NAND3X1 NAND3X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_4917_), .B(_7621_), .C(_5110_), .Y(_5111_) );
OAI21X1 OAI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .B(_5108_), .C(_4842_), .Y(_5112_) );
NAND3X1 NAND3X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_4840_), .B(_5097_), .C(_5101_), .Y(_5113_) );
NAND3X1 NAND3X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_7621_), .B(_5113_), .C(_5112_), .Y(_5114_) );
NAND2X1 NAND2X1_704 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_149_), .B(_5114_), .Y(_5115_) );
NAND3X1 NAND3X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_4916_), .B(_5111_), .C(_5115_), .Y(_5116_) );
NOR2X1 NOR2X1_399 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_149_), .B(_5114_), .Y(_5117_) );
AOI21X1 AOI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(_7621_), .B(_5110_), .C(_4917_), .Y(_5118_) );
OAI21X1 OAI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_5117_), .B(_5118_), .C(_4613_), .Y(_5119_) );
NAND3X1 NAND3X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .B(_4915_), .C(_5119_), .Y(_5120_) );
OAI21X1 OAI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(_4615_), .B(_8193_), .C(_4618_), .Y(_5121_) );
OAI21X1 OAI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_5117_), .B(_5118_), .C(_4916_), .Y(_5122_) );
NAND3X1 NAND3X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_4613_), .B(_5111_), .C(_5115_), .Y(_5123_) );
NAND3X1 NAND3X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .B(_5122_), .C(_5121_), .Y(_5124_) );
NAND3X1 NAND3X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_4914_), .B(_5120_), .C(_5124_), .Y(_5125_) );
AOI21X1 AOI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .B(_5122_), .C(_5121_), .Y(_5126_) );
AOI21X1 AOI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .B(_5119_), .C(_4915_), .Y(_5127_) );
OAI21X1 OAI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_5127_), .C(_4848_), .Y(_5128_) );
NAND2X1 NAND2X1_705 ( .gnd(gnd), .vdd(vdd), .A(_5125_), .B(_5128_), .Y(_5129_) );
NAND3X1 NAND3X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_4913_), .B(_7705_), .C(_5129_), .Y(_5130_) );
OAI21X1 OAI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_5127_), .C(_4914_), .Y(_5131_) );
NAND3X1 NAND3X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_4848_), .B(_5120_), .C(_5124_), .Y(_5132_) );
NAND3X1 NAND3X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_7705_), .B(_5132_), .C(_5131_), .Y(_5133_) );
NAND2X1 NAND2X1_706 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_165_), .B(_5133_), .Y(_5134_) );
NAND3X1 NAND3X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_4912_), .B(_5130_), .C(_5134_), .Y(_5135_) );
NOR2X1 NOR2X1_400 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_165_), .B(_5133_), .Y(_5136_) );
AOI21X1 AOI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_7705_), .B(_5129_), .C(_4913_), .Y(_5137_) );
OAI21X1 OAI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(_5136_), .B(_5137_), .C(_4639_), .Y(_5138_) );
NAND3X1 NAND3X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .B(_5135_), .C(_5138_), .Y(_5139_) );
OAI21X1 OAI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(_8192_), .B(_4641_), .C(_4643_), .Y(_5140_) );
OAI21X1 OAI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(_5136_), .B(_5137_), .C(_4912_), .Y(_5141_) );
NAND3X1 NAND3X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_4639_), .B(_5130_), .C(_5134_), .Y(_5142_) );
NAND3X1 NAND3X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_5142_), .B(_5140_), .C(_5141_), .Y(_5143_) );
NAND3X1 NAND3X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_4856_), .B(_5139_), .C(_5143_), .Y(_5144_) );
NAND2X1 NAND2X1_707 ( .gnd(gnd), .vdd(vdd), .A(_5139_), .B(_5143_), .Y(_5145_) );
AOI21X1 AOI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(_4857_), .B(_5145_), .C(_7714_), .Y(_5146_) );
NAND3X1 NAND3X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .B(_5144_), .C(_5146_), .Y(_5147_) );
AOI21X1 AOI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_5142_), .B(_5141_), .C(_5140_), .Y(_5148_) );
AOI21X1 AOI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_5135_), .B(_5138_), .C(_4911_), .Y(_5149_) );
OAI21X1 OAI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(_5148_), .B(_5149_), .C(_4857_), .Y(_5150_) );
NAND3X1 NAND3X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_7713_), .B(_5144_), .C(_5150_), .Y(_5151_) );
NAND2X1 NAND2X1_708 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_181_), .B(_5151_), .Y(_5152_) );
NAND3X1 NAND3X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_4909_), .B(_5147_), .C(_5152_), .Y(_5153_) );
NOR2X1 NOR2X1_401 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_181_), .B(_5151_), .Y(_5154_) );
AOI21X1 AOI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_5144_), .B(_5146_), .C(_4910_), .Y(_5155_) );
OAI21X1 OAI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(_5154_), .B(_5155_), .C(_4657_), .Y(_5156_) );
NAND3X1 NAND3X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_4908_), .B(_5153_), .C(_5156_), .Y(_5157_) );
OAI21X1 OAI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(_4659_), .B(_8189_), .C(_4662_), .Y(_5158_) );
OAI21X1 OAI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(_5154_), .B(_5155_), .C(_4909_), .Y(_5159_) );
NAND3X1 NAND3X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_4657_), .B(_5147_), .C(_5152_), .Y(_5160_) );
NAND3X1 NAND3X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_5160_), .B(_5158_), .C(_5159_), .Y(_5161_) );
NAND3X1 NAND3X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_4865_), .B(_5157_), .C(_5161_), .Y(_5162_) );
AOI21X1 AOI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(_5160_), .B(_5159_), .C(_5158_), .Y(_5163_) );
AOI21X1 AOI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(_5153_), .B(_5156_), .C(_4908_), .Y(_5164_) );
OAI21X1 OAI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(_5163_), .B(_5164_), .C(_4864_), .Y(_5165_) );
NAND2X1 NAND2X1_709 ( .gnd(gnd), .vdd(vdd), .A(_5162_), .B(_5165_), .Y(_5166_) );
NAND3X1 NAND3X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_4907_), .B(_7722_), .C(_5166_), .Y(_5167_) );
OAI21X1 OAI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(_5163_), .B(_5164_), .C(_4865_), .Y(_5168_) );
NAND3X1 NAND3X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_4864_), .B(_5157_), .C(_5161_), .Y(_5169_) );
NAND3X1 NAND3X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_7722_), .B(_5169_), .C(_5168_), .Y(_5170_) );
NAND2X1 NAND2X1_710 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_197_), .B(_5170_), .Y(_5171_) );
NAND3X1 NAND3X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_4906_), .B(_5167_), .C(_5171_), .Y(_5172_) );
NOR2X1 NOR2X1_402 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_197_), .B(_5170_), .Y(_5173_) );
AOI21X1 AOI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_7722_), .B(_5166_), .C(_4907_), .Y(_5174_) );
OAI21X1 OAI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(_5173_), .B(_5174_), .C(_4683_), .Y(_5175_) );
NAND3X1 NAND3X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_5172_), .B(_4905_), .C(_5175_), .Y(_5176_) );
OAI21X1 OAI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(_4685_), .B(_8187_), .C(_4688_), .Y(_5177_) );
OAI21X1 OAI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(_5173_), .B(_5174_), .C(_4906_), .Y(_5178_) );
NAND3X1 NAND3X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_4683_), .B(_5167_), .C(_5171_), .Y(_5179_) );
NAND3X1 NAND3X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_5179_), .B(_5178_), .C(_5177_), .Y(_5180_) );
NAND3X1 NAND3X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_4873_), .B(_5176_), .C(_5180_), .Y(_5181_) );
AOI21X1 AOI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(_5179_), .B(_5178_), .C(_5177_), .Y(_5182_) );
AOI21X1 AOI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_5172_), .B(_5175_), .C(_4905_), .Y(_5183_) );
OAI21X1 OAI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(_5182_), .B(_5183_), .C(_4872_), .Y(_5184_) );
NAND2X1 NAND2X1_711 ( .gnd(gnd), .vdd(vdd), .A(_5181_), .B(_5184_), .Y(_5185_) );
NAND3X1 NAND3X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_4904_), .B(_7730_), .C(_5185_), .Y(_5186_) );
OAI21X1 OAI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(_5182_), .B(_5183_), .C(_4873_), .Y(_5187_) );
NAND3X1 NAND3X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_4872_), .B(_5176_), .C(_5180_), .Y(_5188_) );
NAND3X1 NAND3X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_7730_), .B(_5188_), .C(_5187_), .Y(_5189_) );
NAND2X1 NAND2X1_712 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_213_), .B(_5189_), .Y(_5190_) );
NAND3X1 NAND3X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .B(_5186_), .C(_5190_), .Y(_5191_) );
NOR2X1 NOR2X1_403 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_213_), .B(_5189_), .Y(_5192_) );
AOI21X1 AOI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(_7730_), .B(_5185_), .C(_4904_), .Y(_5193_) );
OAI21X1 OAI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_5192_), .B(_5193_), .C(_4704_), .Y(_5194_) );
NAND3X1 NAND3X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_5191_), .B(_4902_), .C(_5194_), .Y(_5195_) );
OAI21X1 OAI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_4706_), .B(_8185_), .C(_4710_), .Y(_5196_) );
OAI21X1 OAI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(_5192_), .B(_5193_), .C(_4903_), .Y(_5197_) );
NAND3X1 NAND3X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_4704_), .B(_5186_), .C(_5190_), .Y(_5198_) );
NAND3X1 NAND3X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_5198_), .B(_5196_), .C(_5197_), .Y(_5199_) );
NAND3X1 NAND3X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .B(_5195_), .C(_5199_), .Y(_5200_) );
AOI21X1 AOI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_5198_), .B(_5197_), .C(_5196_), .Y(_5201_) );
AOI21X1 AOI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(_5191_), .B(_5194_), .C(_4902_), .Y(_5202_) );
OAI21X1 OAI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_5202_), .C(_4880_), .Y(_5203_) );
NAND2X1 NAND2X1_713 ( .gnd(gnd), .vdd(vdd), .A(_5200_), .B(_5203_), .Y(_5204_) );
NAND3X1 NAND3X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_4901_), .B(_7739_), .C(_5204_), .Y(_5205_) );
OAI21X1 OAI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_5202_), .C(_4881_), .Y(_5206_) );
NAND3X1 NAND3X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_4880_), .B(_5195_), .C(_5199_), .Y(_5207_) );
NAND3X1 NAND3X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_7739_), .B(_5207_), .C(_5206_), .Y(_5208_) );
NAND2X1 NAND2X1_714 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_229_), .B(_5208_), .Y(_5209_) );
NAND3X1 NAND3X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_4900_), .B(_5205_), .C(_5209_), .Y(_5210_) );
NOR2X1 NOR2X1_404 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_229_), .B(_5208_), .Y(_5211_) );
AOI21X1 AOI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_7739_), .B(_5204_), .C(_4901_), .Y(_5212_) );
OAI21X1 OAI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_5211_), .B(_5212_), .C(_4731_), .Y(_5213_) );
NAND3X1 NAND3X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .B(_5210_), .C(_5213_), .Y(_5214_) );
OAI21X1 OAI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(_8183_), .B(_4733_), .C(_4736_), .Y(_5215_) );
OAI21X1 OAI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_5211_), .B(_5212_), .C(_4900_), .Y(_5216_) );
NAND3X1 NAND3X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_4731_), .B(_5205_), .C(_5209_), .Y(_5217_) );
NAND3X1 NAND3X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_5215_), .B(_5217_), .C(_5216_), .Y(_5218_) );
NAND3X1 NAND3X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_5214_), .C(_5218_), .Y(_5219_) );
NAND2X1 NAND2X1_715 ( .gnd(gnd), .vdd(vdd), .A(_5214_), .B(_5218_), .Y(_5220_) );
AOI21X1 AOI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(_4889_), .B(_5220_), .C(_7936_), .Y(_5221_) );
NAND3X1 NAND3X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_4898_), .B(_5219_), .C(_5221_), .Y(_5222_) );
AOI21X1 AOI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(_5217_), .B(_5216_), .C(_5215_), .Y(_5223_) );
AOI21X1 AOI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_5210_), .B(_5213_), .C(_4899_), .Y(_5224_) );
OAI21X1 OAI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(_5223_), .B(_5224_), .C(_4889_), .Y(_5225_) );
NAND3X1 NAND3X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_7747_), .B(_5219_), .C(_5225_), .Y(_5226_) );
NAND2X1 NAND2X1_716 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_245_), .B(_5226_), .Y(_5227_) );
NAND3X1 NAND3X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_4748_), .B(_5222_), .C(_5227_), .Y(_5228_) );
INVX1 INVX1_696 ( .gnd(gnd), .vdd(vdd), .A(_4748_), .Y(_5229_) );
NOR2X1 NOR2X1_405 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_245_), .B(_5226_), .Y(_5230_) );
AOI21X1 AOI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_5219_), .B(_5221_), .C(_4898_), .Y(_5231_) );
OAI21X1 OAI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(_5230_), .B(_5231_), .C(_5229_), .Y(_5232_) );
NAND3X1 NAND3X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_5228_), .B(_4897_), .C(_5232_), .Y(_5233_) );
AOI21X1 AOI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_4756_), .B(_8181_), .C(_4760_), .Y(_5234_) );
NOR3X1 NOR3X1_141 ( .gnd(gnd), .vdd(vdd), .A(_5229_), .B(_5231_), .C(_5230_), .Y(_5235_) );
AOI21X1 AOI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(_5222_), .B(_5227_), .C(_4748_), .Y(_5236_) );
OAI21X1 OAI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_5235_), .B(_5236_), .C(_5234_), .Y(_5237_) );
NAND3X1 NAND3X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .B(_5233_), .C(_5237_), .Y(_5238_) );
INVX1 INVX1_697 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .Y(_5239_) );
NAND3X1 NAND3X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_5228_), .B(_5234_), .C(_5232_), .Y(_5240_) );
OAI21X1 OAI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(_5235_), .B(_5236_), .C(_4897_), .Y(_5241_) );
NAND3X1 NAND3X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_5239_), .B(_5240_), .C(_5241_), .Y(_5242_) );
NAND2X1 NAND2X1_717 ( .gnd(gnd), .vdd(vdd), .A(_5238_), .B(_5242_), .Y(_5243_) );
XNOR2X1 XNOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_5243_), .B(_4772_), .Y(module_1_H_5_) );
AOI21X1 AOI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_5238_), .B(_5242_), .C(_4772_), .Y(_5244_) );
AOI21X1 AOI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(_5228_), .B(_4897_), .C(_5236_), .Y(_5245_) );
AOI21X1 AOI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_5205_), .B(_5209_), .C(_4731_), .Y(_5246_) );
AOI21X1 AOI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(_5217_), .B(_5215_), .C(_5246_), .Y(_5247_) );
INVX1 INVX1_698 ( .gnd(gnd), .vdd(vdd), .A(_7917_), .Y(_5248_) );
INVX1 INVX1_699 ( .gnd(gnd), .vdd(vdd), .A(_7918_), .Y(_5249_) );
NOR2X1 NOR2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_5249_), .B(_5248_), .Y(_5250_) );
INVX1 INVX1_700 ( .gnd(gnd), .vdd(vdd), .A(_5250_), .Y(_5251_) );
AOI21X1 AOI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_5186_), .B(_5190_), .C(_4704_), .Y(_5252_) );
AOI21X1 AOI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(_5198_), .B(_5196_), .C(_5252_), .Y(_5253_) );
INVX1 INVX1_701 ( .gnd(gnd), .vdd(vdd), .A(_7907_), .Y(_5254_) );
AOI21X1 AOI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_5167_), .B(_5171_), .C(_4683_), .Y(_5255_) );
AOI21X1 AOI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(_5179_), .B(_5177_), .C(_5255_), .Y(_5256_) );
NOR2X1 NOR2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_7897_), .B(_7896_), .Y(_5257_) );
INVX2 INVX2_177 ( .gnd(gnd), .vdd(vdd), .A(_5257_), .Y(_5258_) );
NOR3X1 NOR3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_4909_), .B(_5155_), .C(_5154_), .Y(_5259_) );
OAI21X1 OAI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_5259_), .B(_4908_), .C(_5159_), .Y(_5260_) );
INVX2 INVX2_178 ( .gnd(gnd), .vdd(vdd), .A(_7889_), .Y(_5261_) );
AOI21X1 AOI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_5130_), .B(_5134_), .C(_4639_), .Y(_5262_) );
AOI21X1 AOI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_5142_), .B(_5140_), .C(_5262_), .Y(_5263_) );
INVX1 INVX1_702 ( .gnd(gnd), .vdd(vdd), .A(_5122_), .Y(_5264_) );
AOI21X1 AOI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .B(_5121_), .C(_5264_), .Y(_5265_) );
NOR2X1 NOR2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_7868_), .B(_7869_), .Y(_5266_) );
INVX1 INVX1_703 ( .gnd(gnd), .vdd(vdd), .A(_5266_), .Y(_5267_) );
OAI21X1 OAI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(_5096_), .B(_4918_), .C(_5103_), .Y(_5268_) );
INVX2 INVX2_179 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .Y(_5269_) );
AOI21X1 AOI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_5071_), .B(_5067_), .C(_4562_), .Y(_5270_) );
OAI21X1 OAI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_5270_), .B(_4920_), .C(_5079_), .Y(_5271_) );
INVX2 INVX2_180 ( .gnd(gnd), .vdd(vdd), .A(_5067_), .Y(_5272_) );
NAND2X1 NAND2X1_718 ( .gnd(gnd), .vdd(vdd), .A(_5051_), .B(_5064_), .Y(_5273_) );
INVX2 INVX2_181 ( .gnd(gnd), .vdd(vdd), .A(_5046_), .Y(_5274_) );
NAND2X1 NAND2X1_719 ( .gnd(gnd), .vdd(vdd), .A(_5037_), .B(_5039_), .Y(_5275_) );
INVX2 INVX2_182 ( .gnd(gnd), .vdd(vdd), .A(_5025_), .Y(_5276_) );
NAND2X1 NAND2X1_720 ( .gnd(gnd), .vdd(vdd), .A(_5016_), .B(_5018_), .Y(_5277_) );
INVX2 INVX2_183 ( .gnd(gnd), .vdd(vdd), .A(_5004_), .Y(_5278_) );
NAND2X1 NAND2X1_721 ( .gnd(gnd), .vdd(vdd), .A(_4994_), .B(_4996_), .Y(_5279_) );
INVX2 INVX2_184 ( .gnd(gnd), .vdd(vdd), .A(_4982_), .Y(_5280_) );
INVX1 INVX1_704 ( .gnd(gnd), .vdd(vdd), .A(_4974_), .Y(_5281_) );
OAI21X1 OAI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_5281_), .B(_4930_), .C(_4973_), .Y(_5282_) );
INVX2 INVX2_185 ( .gnd(gnd), .vdd(vdd), .A(_4962_), .Y(_5283_) );
NAND3X1 NAND3X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_8225_), .B(_4942_), .C(_4946_), .Y(_5284_) );
INVX1 INVX1_705 ( .gnd(gnd), .vdd(vdd), .A(_4942_), .Y(_5285_) );
NAND2X1 NAND2X1_722 ( .gnd(gnd), .vdd(vdd), .A(_7764_), .B(_7768_), .Y(_5286_) );
INVX1 INVX1_706 ( .gnd(gnd), .vdd(vdd), .A(_5286_), .Y(_5287_) );
INVX1 INVX1_707 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_6_), .Y(_5288_) );
AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_4939_), .B(_5288_), .Y(_5289_) );
NOR2X1 NOR2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_5288_), .B(_4939_), .Y(_5290_) );
OAI21X1 OAI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(_5289_), .B(_5290_), .C(_5287_), .Y(_5291_) );
NOR2X1 NOR2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_5290_), .B(_5289_), .Y(_5292_) );
OAI21X1 OAI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_7765_), .B(_7766_), .C(_5292_), .Y(_5293_) );
NAND3X1 NAND3X1_1146 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_22_), .B(_5291_), .C(_5293_), .Y(_5294_) );
INVX1 INVX1_708 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_22_), .Y(_5295_) );
OAI21X1 OAI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_5289_), .B(_5290_), .C(_5286_), .Y(_5296_) );
NAND2X1 NAND2X1_723 ( .gnd(gnd), .vdd(vdd), .A(_5287_), .B(_5292_), .Y(_5297_) );
NAND3X1 NAND3X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_5295_), .B(_5296_), .C(_5297_), .Y(_5298_) );
NAND3X1 NAND3X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_5285_), .B(_5298_), .C(_5294_), .Y(_5299_) );
AOI21X1 AOI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_5296_), .B(_5297_), .C(_5295_), .Y(_5300_) );
AOI21X1 AOI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_5291_), .B(_5293_), .C(module_1_W_22_), .Y(_5301_) );
OAI21X1 OAI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(_5301_), .B(_5300_), .C(_4942_), .Y(_5302_) );
NAND2X1 NAND2X1_724 ( .gnd(gnd), .vdd(vdd), .A(_5299_), .B(_5302_), .Y(_5303_) );
AOI21X1 AOI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_5284_), .B(_4954_), .C(_5303_), .Y(_5304_) );
INVX1 INVX1_709 ( .gnd(gnd), .vdd(vdd), .A(_5304_), .Y(_5305_) );
OAI21X1 OAI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(_4932_), .B(_4951_), .C(_5284_), .Y(_5306_) );
INVX1 INVX1_710 ( .gnd(gnd), .vdd(vdd), .A(_5303_), .Y(_5307_) );
OR2X2 OR2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_5307_), .B(_5306_), .Y(_5308_) );
INVX2 INVX2_186 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_10_), .Y(_5309_) );
NOR2X1 NOR2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_7777_), .B(_7775_), .Y(_5310_) );
XNOR2X1 XNOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_5310_), .B(_5309_), .Y(_5311_) );
NAND3X1 NAND3X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_5305_), .B(_5311_), .C(_5308_), .Y(_5312_) );
NOR2X1 NOR2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_5306_), .B(_5307_), .Y(_5313_) );
INVX1 INVX1_711 ( .gnd(gnd), .vdd(vdd), .A(_5311_), .Y(_5314_) );
OAI21X1 OAI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(_5313_), .B(_5304_), .C(_5314_), .Y(_5315_) );
NAND3X1 NAND3X1_1150 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf3_), .B(_5315_), .C(_5312_), .Y(_5316_) );
INVX2 INVX2_187 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf2_), .Y(_5317_) );
NAND3X1 NAND3X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_5305_), .B(_5314_), .C(_5308_), .Y(_5318_) );
OAI21X1 OAI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_5313_), .B(_5304_), .C(_5311_), .Y(_5319_) );
NAND3X1 NAND3X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_5317_), .B(_5319_), .C(_5318_), .Y(_5320_) );
NAND3X1 NAND3X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_5283_), .B(_5316_), .C(_5320_), .Y(_5321_) );
NAND3X1 NAND3X1_1154 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf1_), .B(_5319_), .C(_5318_), .Y(_5322_) );
NAND3X1 NAND3X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_5317_), .B(_5315_), .C(_5312_), .Y(_5323_) );
NAND3X1 NAND3X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_4962_), .B(_5322_), .C(_5323_), .Y(_5324_) );
NAND3X1 NAND3X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_5282_), .B(_5321_), .C(_5324_), .Y(_5325_) );
INVX1 INVX1_712 ( .gnd(gnd), .vdd(vdd), .A(_4973_), .Y(_5326_) );
NOR2X1 NOR2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_5326_), .B(_4980_), .Y(_5327_) );
AOI21X1 AOI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_5322_), .B(_5323_), .C(_4962_), .Y(_5328_) );
AOI21X1 AOI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_5316_), .B(_5320_), .C(_5283_), .Y(_5329_) );
OAI21X1 OAI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_5328_), .B(_5329_), .C(_5327_), .Y(_5330_) );
NOR2X1 NOR2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_7787_), .B(_7794_), .Y(_5331_) );
NAND2X1 NAND2X1_725 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_26_), .B(module_1_W_10_), .Y(_5332_) );
INVX1 INVX1_713 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_26_), .Y(_5333_) );
NAND2X1 NAND2X1_726 ( .gnd(gnd), .vdd(vdd), .A(_5333_), .B(_5309_), .Y(_5334_) );
AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_5334_), .B(_5332_), .Y(_5335_) );
NAND2X1 NAND2X1_727 ( .gnd(gnd), .vdd(vdd), .A(_4792_), .B(_5335_), .Y(_5336_) );
NAND2X1 NAND2X1_728 ( .gnd(gnd), .vdd(vdd), .A(_5332_), .B(_5334_), .Y(_5337_) );
OAI21X1 OAI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(_4790_), .B(_4791_), .C(_5337_), .Y(_5338_) );
NAND3X1 NAND3X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_5336_), .B(_5338_), .C(_4796_), .Y(_5339_) );
OAI21X1 OAI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_24_), .B(module_1_W_8_), .C(_4794_), .Y(_5340_) );
INVX1 INVX1_714 ( .gnd(gnd), .vdd(vdd), .A(_4792_), .Y(_5341_) );
NOR2X1 NOR2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_5341_), .B(_5337_), .Y(_5342_) );
NOR2X1 NOR2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_4792_), .B(_5335_), .Y(_5343_) );
OAI21X1 OAI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(_5343_), .B(_5342_), .C(_5340_), .Y(_5344_) );
NAND2X1 NAND2X1_729 ( .gnd(gnd), .vdd(vdd), .A(_5344_), .B(_5339_), .Y(_5345_) );
XNOR2X1 XNOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_5331_), .B(_5345_), .Y(_5346_) );
NAND3X1 NAND3X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_5325_), .B(_5346_), .C(_5330_), .Y(_5347_) );
NAND3X1 NAND3X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_4962_), .B(_5316_), .C(_5320_), .Y(_5348_) );
NAND3X1 NAND3X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_5283_), .B(_5322_), .C(_5323_), .Y(_5349_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_4973_), .B(_4975_), .C(_5348_), .D(_5349_), .Y(_5350_) );
AOI21X1 AOI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_5321_), .B(_5324_), .C(_5282_), .Y(_5351_) );
INVX1 INVX1_715 ( .gnd(gnd), .vdd(vdd), .A(_5346_), .Y(_5352_) );
OAI21X1 OAI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(_5350_), .B(_5351_), .C(_5352_), .Y(_5353_) );
NAND3X1 NAND3X1_1162 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf3_), .B(_5347_), .C(_5353_), .Y(_5354_) );
INVX1 INVX1_716 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf2_), .Y(_5355_) );
NAND3X1 NAND3X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_5325_), .B(_5352_), .C(_5330_), .Y(_5356_) );
OAI21X1 OAI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_5350_), .B(_5351_), .C(_5346_), .Y(_5357_) );
NAND3X1 NAND3X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_5355_), .B(_5356_), .C(_5357_), .Y(_5358_) );
NAND3X1 NAND3X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_5280_), .B(_5354_), .C(_5358_), .Y(_5359_) );
NAND3X1 NAND3X1_1166 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf1_), .B(_5356_), .C(_5357_), .Y(_5360_) );
NAND3X1 NAND3X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_5355_), .B(_5347_), .C(_5353_), .Y(_5361_) );
NAND3X1 NAND3X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_4982_), .B(_5360_), .C(_5361_), .Y(_5362_) );
NAND3X1 NAND3X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_5359_), .B(_5362_), .C(_5279_), .Y(_5363_) );
AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_4996_), .B(_4994_), .Y(_5364_) );
AOI21X1 AOI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_5360_), .B(_5361_), .C(_4982_), .Y(_5365_) );
AOI21X1 AOI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_5354_), .B(_5358_), .C(_5280_), .Y(_5366_) );
OAI21X1 OAI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_5365_), .B(_5366_), .C(_5364_), .Y(_5367_) );
NOR2X1 NOR2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_7804_), .B(_7801_), .Y(_5368_) );
NOR2X1 NOR2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_4789_), .B(_4803_), .Y(_5369_) );
INVX1 INVX1_717 ( .gnd(gnd), .vdd(vdd), .A(_4801_), .Y(_5370_) );
INVX1 INVX1_718 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .Y(_5371_) );
NAND2X1 NAND2X1_730 ( .gnd(gnd), .vdd(vdd), .A(_5371_), .B(_5345_), .Y(_5372_) );
NAND3X1 NAND3X1_1170 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .B(_5344_), .C(_5339_), .Y(_5373_) );
NAND2X1 NAND2X1_731 ( .gnd(gnd), .vdd(vdd), .A(_5373_), .B(_5372_), .Y(_5374_) );
NOR2X1 NOR2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_5370_), .B(_5374_), .Y(_5375_) );
AOI21X1 AOI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(_5373_), .B(_5372_), .C(_4801_), .Y(_5376_) );
NOR2X1 NOR2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_5376_), .B(_5375_), .Y(_5377_) );
NAND2X1 NAND2X1_732 ( .gnd(gnd), .vdd(vdd), .A(_5369_), .B(_5377_), .Y(_5378_) );
OAI21X1 OAI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_5375_), .B(_5376_), .C(_4804_), .Y(_5379_) );
NAND2X1 NAND2X1_733 ( .gnd(gnd), .vdd(vdd), .A(_5379_), .B(_5378_), .Y(_5380_) );
XNOR2X1 XNOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_5368_), .B(_5380_), .Y(_5381_) );
NAND3X1 NAND3X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_5363_), .B(_5381_), .C(_5367_), .Y(_5382_) );
NAND3X1 NAND3X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_4982_), .B(_5354_), .C(_5358_), .Y(_5383_) );
NAND3X1 NAND3X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_5280_), .B(_5360_), .C(_5361_), .Y(_5384_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_4994_), .B(_4996_), .C(_5383_), .D(_5384_), .Y(_5385_) );
AOI21X1 AOI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(_5359_), .B(_5362_), .C(_5279_), .Y(_5386_) );
INVX1 INVX1_719 ( .gnd(gnd), .vdd(vdd), .A(_5381_), .Y(_5387_) );
OAI21X1 OAI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_5385_), .B(_5386_), .C(_5387_), .Y(_5388_) );
NAND3X1 NAND3X1_1174 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf2_), .B(_5388_), .C(_5382_), .Y(_5389_) );
INVX1 INVX1_720 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf1_), .Y(_5390_) );
NAND3X1 NAND3X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_5363_), .B(_5387_), .C(_5367_), .Y(_5391_) );
OAI21X1 OAI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_5385_), .B(_5386_), .C(_5381_), .Y(_5392_) );
NAND3X1 NAND3X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_5390_), .B(_5392_), .C(_5391_), .Y(_5393_) );
NAND3X1 NAND3X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_5278_), .B(_5389_), .C(_5393_), .Y(_5394_) );
NAND3X1 NAND3X1_1178 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf0_), .B(_5392_), .C(_5391_), .Y(_5395_) );
NAND3X1 NAND3X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_5390_), .B(_5388_), .C(_5382_), .Y(_5396_) );
NAND3X1 NAND3X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_5004_), .B(_5395_), .C(_5396_), .Y(_5397_) );
NAND3X1 NAND3X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_5394_), .B(_5397_), .C(_5277_), .Y(_5398_) );
AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_5018_), .B(_5016_), .Y(_5399_) );
AOI21X1 AOI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_5395_), .B(_5396_), .C(_5004_), .Y(_5400_) );
AOI21X1 AOI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_5389_), .B(_5393_), .C(_5278_), .Y(_5401_) );
OAI21X1 OAI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_5400_), .B(_5401_), .C(_5399_), .Y(_5402_) );
INVX2 INVX2_188 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf3_), .Y(_5403_) );
AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_5377_), .B(_5369_), .Y(_5404_) );
INVX1 INVX1_721 ( .gnd(gnd), .vdd(vdd), .A(_5379_), .Y(_5405_) );
OAI21X1 OAI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_5404_), .B(_5405_), .C(_5403_), .Y(_5406_) );
OR2X2 OR2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_5380_), .B(_5403_), .Y(_5407_) );
NAND3X1 NAND3X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_4807_), .B(_5406_), .C(_5407_), .Y(_5408_) );
INVX1 INVX1_722 ( .gnd(gnd), .vdd(vdd), .A(_4807_), .Y(_5409_) );
INVX1 INVX1_723 ( .gnd(gnd), .vdd(vdd), .A(_5406_), .Y(_5410_) );
NOR2X1 NOR2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_5403_), .B(_5380_), .Y(_5411_) );
OAI21X1 OAI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_5410_), .B(_5411_), .C(_5409_), .Y(_5412_) );
NAND2X1 NAND2X1_734 ( .gnd(gnd), .vdd(vdd), .A(_5408_), .B(_5412_), .Y(_5413_) );
OR2X2 OR2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_5413_), .B(_4810_), .Y(_5414_) );
NOR3X1 NOR3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_5409_), .B(_5411_), .C(_5410_), .Y(_5415_) );
AOI21X1 AOI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(_5406_), .B(_5407_), .C(_4807_), .Y(_5416_) );
OAI21X1 OAI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(_5415_), .B(_5416_), .C(_4810_), .Y(_5417_) );
NAND2X1 NAND2X1_735 ( .gnd(gnd), .vdd(vdd), .A(_5417_), .B(_5414_), .Y(_5418_) );
XNOR2X1 XNOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_8033_), .B(_5418_), .Y(_5419_) );
NAND3X1 NAND3X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_5398_), .B(_5419_), .C(_5402_), .Y(_5420_) );
NAND3X1 NAND3X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_5004_), .B(_5389_), .C(_5393_), .Y(_5421_) );
NAND3X1 NAND3X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_5278_), .B(_5395_), .C(_5396_), .Y(_5422_) );
AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_5016_), .B(_5018_), .C(_5421_), .D(_5422_), .Y(_5423_) );
AOI21X1 AOI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_5394_), .B(_5397_), .C(_5277_), .Y(_5424_) );
INVX1 INVX1_724 ( .gnd(gnd), .vdd(vdd), .A(_5419_), .Y(_5425_) );
OAI21X1 OAI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_5423_), .B(_5424_), .C(_5425_), .Y(_5426_) );
NAND3X1 NAND3X1_1186 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf2_), .B(_5420_), .C(_5426_), .Y(_5427_) );
INVX1 INVX1_725 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf1_), .Y(_5428_) );
OAI21X1 OAI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_5423_), .B(_5424_), .C(_5419_), .Y(_5429_) );
NAND3X1 NAND3X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_5398_), .B(_5425_), .C(_5402_), .Y(_5430_) );
NAND3X1 NAND3X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_5428_), .B(_5430_), .C(_5429_), .Y(_5431_) );
NAND3X1 NAND3X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_5276_), .B(_5427_), .C(_5431_), .Y(_5432_) );
NAND3X1 NAND3X1_1190 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf0_), .B(_5430_), .C(_5429_), .Y(_5433_) );
NAND3X1 NAND3X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_5428_), .B(_5420_), .C(_5426_), .Y(_5434_) );
NAND3X1 NAND3X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_5025_), .B(_5433_), .C(_5434_), .Y(_5435_) );
NAND3X1 NAND3X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_5432_), .B(_5435_), .C(_5275_), .Y(_5436_) );
AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_5039_), .B(_5037_), .Y(_5437_) );
AOI21X1 AOI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_5433_), .B(_5434_), .C(_5025_), .Y(_5438_) );
AOI21X1 AOI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(_5427_), .B(_5431_), .C(_5276_), .Y(_5439_) );
OAI21X1 OAI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_5438_), .B(_5439_), .C(_5437_), .Y(_5440_) );
INVX1 INVX1_726 ( .gnd(gnd), .vdd(vdd), .A(_4815_), .Y(_5441_) );
INVX1 INVX1_727 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf2_), .Y(_5442_) );
NOR2X1 NOR2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_4810_), .B(_5413_), .Y(_5443_) );
INVX1 INVX1_728 ( .gnd(gnd), .vdd(vdd), .A(_5417_), .Y(_5444_) );
OAI21X1 OAI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(_5444_), .B(_5443_), .C(_5442_), .Y(_5445_) );
INVX1 INVX1_729 ( .gnd(gnd), .vdd(vdd), .A(_5445_), .Y(_5446_) );
NOR2X1 NOR2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_5442_), .B(_5418_), .Y(_5447_) );
NOR3X1 NOR3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_5446_), .B(_5441_), .C(_5447_), .Y(_5448_) );
NOR2X1 NOR2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_5443_), .B(_5444_), .Y(_5449_) );
NAND2X1 NAND2X1_736 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf1_), .B(_5449_), .Y(_5450_) );
AOI21X1 AOI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_5445_), .B(_5450_), .C(_4815_), .Y(_5451_) );
NOR3X1 NOR3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_4818_), .B(_5451_), .C(_5448_), .Y(_5452_) );
INVX2 INVX2_189 ( .gnd(gnd), .vdd(vdd), .A(_4818_), .Y(_5453_) );
NAND3X1 NAND3X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_4815_), .B(_5445_), .C(_5450_), .Y(_5454_) );
OAI21X1 OAI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(_5447_), .B(_5446_), .C(_5441_), .Y(_5455_) );
AOI21X1 AOI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(_5454_), .B(_5455_), .C(_5453_), .Y(_5456_) );
NOR2X1 NOR2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_5456_), .B(_5452_), .Y(_5457_) );
OAI21X1 OAI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_7824_), .B(_7825_), .C(_5457_), .Y(_5458_) );
NOR2X1 NOR2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_7825_), .B(_7824_), .Y(_5459_) );
OAI21X1 OAI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(_5452_), .B(_5456_), .C(_5459_), .Y(_5460_) );
NAND2X1 NAND2X1_737 ( .gnd(gnd), .vdd(vdd), .A(_5458_), .B(_5460_), .Y(_5461_) );
NAND3X1 NAND3X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_5436_), .B(_5461_), .C(_5440_), .Y(_5462_) );
NAND3X1 NAND3X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_5025_), .B(_5427_), .C(_5431_), .Y(_5463_) );
NAND3X1 NAND3X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_5276_), .B(_5433_), .C(_5434_), .Y(_5464_) );
AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_5037_), .B(_5039_), .C(_5463_), .D(_5464_), .Y(_5465_) );
AOI21X1 AOI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_5432_), .B(_5435_), .C(_5275_), .Y(_5466_) );
INVX1 INVX1_730 ( .gnd(gnd), .vdd(vdd), .A(_5461_), .Y(_5467_) );
OAI21X1 OAI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(_5465_), .B(_5466_), .C(_5467_), .Y(_5468_) );
NAND3X1 NAND3X1_1198 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf2_), .B(_5462_), .C(_5468_), .Y(_5469_) );
INVX1 INVX1_731 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf1_), .Y(_5470_) );
OAI21X1 OAI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_5465_), .B(_5466_), .C(_5461_), .Y(_5471_) );
NAND3X1 NAND3X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_5436_), .B(_5467_), .C(_5440_), .Y(_5472_) );
NAND3X1 NAND3X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_5470_), .B(_5472_), .C(_5471_), .Y(_5473_) );
NAND3X1 NAND3X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_5274_), .B(_5469_), .C(_5473_), .Y(_5474_) );
NAND3X1 NAND3X1_1202 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf0_), .B(_5472_), .C(_5471_), .Y(_5475_) );
NAND3X1 NAND3X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_5470_), .B(_5462_), .C(_5468_), .Y(_5476_) );
NAND3X1 NAND3X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_5046_), .B(_5475_), .C(_5476_), .Y(_5477_) );
NAND3X1 NAND3X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_5474_), .B(_5477_), .C(_5273_), .Y(_5478_) );
AND2X2 AND2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_5064_), .B(_5051_), .Y(_5479_) );
AOI21X1 AOI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(_5475_), .B(_5476_), .C(_5046_), .Y(_5480_) );
AOI21X1 AOI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(_5469_), .B(_5473_), .C(_5274_), .Y(_5481_) );
OAI21X1 OAI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_5480_), .B(_5481_), .C(_5479_), .Y(_5482_) );
INVX1 INVX1_732 ( .gnd(gnd), .vdd(vdd), .A(_4823_), .Y(_5483_) );
NAND3X1 NAND3X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_5454_), .B(_5455_), .C(_5453_), .Y(_5484_) );
OAI21X1 OAI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_5448_), .B(_5451_), .C(_4818_), .Y(_5485_) );
AOI21X1 AOI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(_5484_), .B(_5485_), .C(bloque_datos_58_bF_buf3_), .Y(_5486_) );
INVX1 INVX1_733 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf2_), .Y(_5487_) );
NOR3X1 NOR3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_5487_), .B(_5456_), .C(_5452_), .Y(_5488_) );
NOR3X1 NOR3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_5483_), .B(_5486_), .C(_5488_), .Y(_5489_) );
OAI21X1 OAI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(_5452_), .B(_5456_), .C(_5487_), .Y(_5490_) );
NAND3X1 NAND3X1_1207 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf1_), .B(_5484_), .C(_5485_), .Y(_5491_) );
AOI21X1 AOI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_5491_), .B(_5490_), .C(_4823_), .Y(_5492_) );
NOR3X1 NOR3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_4826_), .B(_5492_), .C(_5489_), .Y(_5493_) );
NOR2X1 NOR2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_4786_), .B(_4825_), .Y(_5494_) );
NAND3X1 NAND3X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_4823_), .B(_5491_), .C(_5490_), .Y(_5495_) );
OAI21X1 OAI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(_5488_), .B(_5486_), .C(_5483_), .Y(_5496_) );
AOI21X1 AOI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_5495_), .B(_5496_), .C(_5494_), .Y(_5497_) );
NOR2X1 NOR2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_5497_), .B(_5493_), .Y(_5498_) );
OAI21X1 OAI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(_7844_), .B(_7845_), .C(_5498_), .Y(_5499_) );
NOR2X1 NOR2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_7845_), .B(_7844_), .Y(_5500_) );
OAI21X1 OAI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(_5493_), .B(_5497_), .C(_5500_), .Y(_5501_) );
NAND2X1 NAND2X1_738 ( .gnd(gnd), .vdd(vdd), .A(_5499_), .B(_5501_), .Y(_5502_) );
NAND3X1 NAND3X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_5478_), .B(_5502_), .C(_5482_), .Y(_5503_) );
NAND3X1 NAND3X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_5046_), .B(_5469_), .C(_5473_), .Y(_5504_) );
NAND3X1 NAND3X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_5274_), .B(_5475_), .C(_5476_), .Y(_5505_) );
AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_5051_), .B(_5064_), .C(_5504_), .D(_5505_), .Y(_5506_) );
AOI21X1 AOI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(_5474_), .B(_5477_), .C(_5273_), .Y(_5507_) );
INVX1 INVX1_734 ( .gnd(gnd), .vdd(vdd), .A(_5502_), .Y(_5508_) );
OAI21X1 OAI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_5507_), .B(_5506_), .C(_5508_), .Y(_5509_) );
NAND3X1 NAND3X1_1212 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf3_), .B(_5509_), .C(_5503_), .Y(_5510_) );
INVX1 INVX1_735 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf2_), .Y(_5511_) );
OAI21X1 OAI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_5507_), .B(_5506_), .C(_5502_), .Y(_5512_) );
NAND3X1 NAND3X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_5478_), .B(_5508_), .C(_5482_), .Y(_5513_) );
NAND3X1 NAND3X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_5511_), .B(_5512_), .C(_5513_), .Y(_5514_) );
NAND3X1 NAND3X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_5272_), .B(_5510_), .C(_5514_), .Y(_5515_) );
NAND3X1 NAND3X1_1216 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf1_), .B(_5512_), .C(_5513_), .Y(_5516_) );
NAND3X1 NAND3X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_5511_), .B(_5509_), .C(_5503_), .Y(_5517_) );
NAND3X1 NAND3X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_5067_), .B(_5516_), .C(_5517_), .Y(_5518_) );
NAND3X1 NAND3X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_5271_), .B(_5515_), .C(_5518_), .Y(_5519_) );
INVX1 INVX1_736 ( .gnd(gnd), .vdd(vdd), .A(_5271_), .Y(_5520_) );
AOI21X1 AOI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(_5516_), .B(_5517_), .C(_5067_), .Y(_5521_) );
AOI21X1 AOI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_5510_), .B(_5514_), .C(_5272_), .Y(_5522_) );
OAI21X1 OAI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_5521_), .B(_5522_), .C(_5520_), .Y(_5523_) );
INVX1 INVX1_737 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf3_), .Y(_5524_) );
OAI21X1 OAI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_5493_), .B(_5497_), .C(_5524_), .Y(_5525_) );
NAND3X1 NAND3X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_5494_), .B(_5495_), .C(_5496_), .Y(_5526_) );
OAI21X1 OAI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_5489_), .B(_5492_), .C(_4826_), .Y(_5527_) );
NAND3X1 NAND3X1_1221 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf2_), .B(_5526_), .C(_5527_), .Y(_5528_) );
NAND2X1 NAND2X1_739 ( .gnd(gnd), .vdd(vdd), .A(_5528_), .B(_5525_), .Y(_5529_) );
NOR2X1 NOR2X1_430 ( .gnd(gnd), .vdd(vdd), .A(_4829_), .B(_5529_), .Y(_5530_) );
INVX1 INVX1_738 ( .gnd(gnd), .vdd(vdd), .A(_4829_), .Y(_5531_) );
AOI21X1 AOI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(_5528_), .B(_5525_), .C(_5531_), .Y(_5532_) );
NOR3X1 NOR3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_4832_), .B(_5532_), .C(_5530_), .Y(_5533_) );
NOR2X1 NOR2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_4570_), .B(_4830_), .Y(_5534_) );
NAND3X1 NAND3X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_5525_), .B(_5528_), .C(_5531_), .Y(_5535_) );
INVX1 INVX1_739 ( .gnd(gnd), .vdd(vdd), .A(_5532_), .Y(_5536_) );
AOI21X1 AOI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_5535_), .B(_5536_), .C(_5534_), .Y(_5537_) );
NOR2X1 NOR2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_5537_), .B(_5533_), .Y(_5538_) );
OAI21X1 OAI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_7856_), .B(_7857_), .C(_5538_), .Y(_5539_) );
NOR2X1 NOR2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_7857_), .B(_7856_), .Y(_5540_) );
OAI21X1 OAI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(_5533_), .B(_5537_), .C(_5540_), .Y(_5541_) );
NAND2X1 NAND2X1_740 ( .gnd(gnd), .vdd(vdd), .A(_5539_), .B(_5541_), .Y(_5542_) );
NAND3X1 NAND3X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_5519_), .B(_5542_), .C(_5523_), .Y(_5543_) );
NAND3X1 NAND3X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_5067_), .B(_5510_), .C(_5514_), .Y(_5544_) );
NAND3X1 NAND3X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_5272_), .B(_5516_), .C(_5517_), .Y(_5545_) );
AOI21X1 AOI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(_5544_), .B(_5545_), .C(_5520_), .Y(_5546_) );
AOI21X1 AOI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(_5515_), .B(_5518_), .C(_5271_), .Y(_5547_) );
INVX1 INVX1_740 ( .gnd(gnd), .vdd(vdd), .A(_5542_), .Y(_5548_) );
OAI21X1 OAI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_5547_), .C(_5548_), .Y(_5549_) );
NAND3X1 NAND3X1_1226 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_134_), .B(_5543_), .C(_5549_), .Y(_5550_) );
INVX1 INVX1_741 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_134_), .Y(_5551_) );
NAND3X1 NAND3X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_5519_), .B(_5548_), .C(_5523_), .Y(_5552_) );
OAI21X1 OAI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_5547_), .C(_5542_), .Y(_5553_) );
NAND3X1 NAND3X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_5551_), .B(_5552_), .C(_5553_), .Y(_5554_) );
NAND3X1 NAND3X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_5269_), .B(_5550_), .C(_5554_), .Y(_5555_) );
NAND3X1 NAND3X1_1230 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_134_), .B(_5552_), .C(_5553_), .Y(_5556_) );
NAND3X1 NAND3X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_5551_), .B(_5543_), .C(_5549_), .Y(_5557_) );
NAND3X1 NAND3X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_5556_), .C(_5557_), .Y(_5558_) );
NAND3X1 NAND3X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_5268_), .B(_5555_), .C(_5558_), .Y(_5559_) );
INVX2 INVX2_190 ( .gnd(gnd), .vdd(vdd), .A(_5268_), .Y(_5560_) );
AOI21X1 AOI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(_5556_), .B(_5557_), .C(_5094_), .Y(_5561_) );
AOI21X1 AOI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(_5550_), .B(_5554_), .C(_5269_), .Y(_5562_) );
OAI21X1 OAI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(_5561_), .B(_5562_), .C(_5560_), .Y(_5563_) );
INVX1 INVX1_742 ( .gnd(gnd), .vdd(vdd), .A(_4835_), .Y(_5564_) );
INVX1 INVX1_743 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf2_), .Y(_5565_) );
OAI21X1 OAI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_5533_), .B(_5537_), .C(_5565_), .Y(_5566_) );
NAND3X1 NAND3X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_5534_), .B(_5535_), .C(_5536_), .Y(_5567_) );
OAI21X1 OAI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_5530_), .B(_5532_), .C(_4832_), .Y(_5568_) );
NAND3X1 NAND3X1_1235 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf1_), .B(_5568_), .C(_5567_), .Y(_5569_) );
NAND3X1 NAND3X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_5566_), .B(_5569_), .C(_5564_), .Y(_5570_) );
AOI21X1 AOI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(_5568_), .B(_5567_), .C(bloque_datos_90_bF_buf0_), .Y(_5571_) );
NOR3X1 NOR3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_5537_), .B(_5565_), .C(_5533_), .Y(_5572_) );
OAI21X1 OAI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(_5572_), .B(_5571_), .C(_4835_), .Y(_5573_) );
AND2X2 AND2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_5573_), .B(_5570_), .Y(_5574_) );
NAND2X1 NAND2X1_741 ( .gnd(gnd), .vdd(vdd), .A(_4838_), .B(_5574_), .Y(_5575_) );
INVX1 INVX1_744 ( .gnd(gnd), .vdd(vdd), .A(_5575_), .Y(_5576_) );
NOR2X1 NOR2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_4838_), .B(_5574_), .Y(_5577_) );
NOR2X1 NOR2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_5577_), .B(_5576_), .Y(_5578_) );
INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(_5578_), .Y(_5579_) );
NAND3X1 NAND3X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_5559_), .B(_5579_), .C(_5563_), .Y(_5580_) );
NAND3X1 NAND3X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_5550_), .C(_5554_), .Y(_5581_) );
NAND3X1 NAND3X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_5269_), .B(_5556_), .C(_5557_), .Y(_5582_) );
AOI21X1 AOI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(_5581_), .B(_5582_), .C(_5560_), .Y(_5583_) );
AOI21X1 AOI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(_5555_), .B(_5558_), .C(_5268_), .Y(_5584_) );
OAI21X1 OAI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(_5583_), .B(_5584_), .C(_5578_), .Y(_5585_) );
NAND3X1 NAND3X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_5267_), .B(_5580_), .C(_5585_), .Y(_5586_) );
NAND2X1 NAND2X1_742 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_150_), .B(_5586_), .Y(_5587_) );
INVX2 INVX2_191 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_150_), .Y(_5588_) );
OAI21X1 OAI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(_5583_), .B(_5584_), .C(_5579_), .Y(_5589_) );
NAND3X1 NAND3X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_5559_), .B(_5578_), .C(_5563_), .Y(_5590_) );
AOI21X1 AOI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(_5590_), .B(_5589_), .C(_5266_), .Y(_5591_) );
NAND2X1 NAND2X1_743 ( .gnd(gnd), .vdd(vdd), .A(_5588_), .B(_5591_), .Y(_5592_) );
NAND3X1 NAND3X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_5117_), .B(_5587_), .C(_5592_), .Y(_5593_) );
NAND2X1 NAND2X1_744 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_150_), .B(_5591_), .Y(_5594_) );
NAND2X1 NAND2X1_745 ( .gnd(gnd), .vdd(vdd), .A(_5588_), .B(_5586_), .Y(_5595_) );
NAND3X1 NAND3X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_5111_), .B(_5595_), .C(_5594_), .Y(_5596_) );
AOI21X1 AOI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(_5593_), .B(_5596_), .C(_5265_), .Y(_5597_) );
INVX1 INVX1_745 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .Y(_5598_) );
OAI21X1 OAI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(_5598_), .B(_4915_), .C(_5122_), .Y(_5599_) );
NAND3X1 NAND3X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_5111_), .B(_5587_), .C(_5592_), .Y(_5600_) );
NAND3X1 NAND3X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_5117_), .B(_5595_), .C(_5594_), .Y(_5601_) );
AOI21X1 AOI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(_5600_), .B(_5601_), .C(_5599_), .Y(_5602_) );
INVX1 INVX1_746 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_138_), .Y(_5603_) );
OAI21X1 OAI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(_5576_), .B(_5577_), .C(_5603_), .Y(_5604_) );
NAND2X1 NAND2X1_746 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_138_), .B(_5578_), .Y(_5605_) );
NAND2X1 NAND2X1_747 ( .gnd(gnd), .vdd(vdd), .A(_5604_), .B(_5605_), .Y(_5606_) );
NOR2X1 NOR2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_4843_), .B(_5606_), .Y(_5607_) );
INVX1 INVX1_747 ( .gnd(gnd), .vdd(vdd), .A(_5607_), .Y(_5608_) );
OAI21X1 OAI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(_4781_), .B(_4840_), .C(_5606_), .Y(_5609_) );
NAND3X1 NAND3X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_4846_), .B(_5609_), .C(_5608_), .Y(_5610_) );
INVX1 INVX1_748 ( .gnd(gnd), .vdd(vdd), .A(_5609_), .Y(_5611_) );
OAI21X1 OAI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(_5611_), .B(_5607_), .C(_4847_), .Y(_5612_) );
NAND2X1 NAND2X1_748 ( .gnd(gnd), .vdd(vdd), .A(_5612_), .B(_5610_), .Y(_5613_) );
INVX2 INVX2_192 ( .gnd(gnd), .vdd(vdd), .A(_5613_), .Y(_5614_) );
OAI21X1 OAI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(_5597_), .B(_5602_), .C(_5614_), .Y(_5615_) );
NAND3X1 NAND3X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_5600_), .B(_5601_), .C(_5599_), .Y(_5616_) );
AOI21X1 AOI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(_5595_), .B(_5594_), .C(_5117_), .Y(_5617_) );
AOI21X1 AOI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(_5587_), .B(_5592_), .C(_5111_), .Y(_5618_) );
OAI21X1 OAI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(_5617_), .B(_5618_), .C(_5265_), .Y(_5619_) );
NAND3X1 NAND3X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_5613_), .B(_5616_), .C(_5619_), .Y(_5620_) );
NAND3X1 NAND3X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_8092_), .B(_5620_), .C(_5615_), .Y(_5621_) );
NAND2X1 NAND2X1_749 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_166_), .B(_5621_), .Y(_5622_) );
INVX2 INVX2_193 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_166_), .Y(_5623_) );
NAND3X1 NAND3X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_5614_), .B(_5616_), .C(_5619_), .Y(_5624_) );
OAI21X1 OAI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(_5597_), .B(_5602_), .C(_5613_), .Y(_5625_) );
AOI21X1 AOI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(_5624_), .B(_5625_), .C(_7879_), .Y(_5626_) );
NAND2X1 NAND2X1_750 ( .gnd(gnd), .vdd(vdd), .A(_5623_), .B(_5626_), .Y(_5627_) );
NAND3X1 NAND3X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_5136_), .B(_5622_), .C(_5627_), .Y(_5628_) );
NAND2X1 NAND2X1_751 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_166_), .B(_5626_), .Y(_5629_) );
NAND2X1 NAND2X1_752 ( .gnd(gnd), .vdd(vdd), .A(_5623_), .B(_5621_), .Y(_5630_) );
NAND3X1 NAND3X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_5130_), .B(_5630_), .C(_5629_), .Y(_5631_) );
AOI21X1 AOI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(_5628_), .B(_5631_), .C(_5263_), .Y(_5632_) );
NOR3X1 NOR3X1_151 ( .gnd(gnd), .vdd(vdd), .A(_5137_), .B(_4912_), .C(_5136_), .Y(_5633_) );
OAI21X1 OAI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(_5633_), .B(_4911_), .C(_5141_), .Y(_5634_) );
NAND3X1 NAND3X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_5130_), .B(_5622_), .C(_5627_), .Y(_5635_) );
NAND3X1 NAND3X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_5136_), .B(_5630_), .C(_5629_), .Y(_5636_) );
AOI21X1 AOI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(_5635_), .B(_5636_), .C(_5634_), .Y(_5637_) );
INVX1 INVX1_749 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_154_), .Y(_5638_) );
NAND2X1 NAND2X1_753 ( .gnd(gnd), .vdd(vdd), .A(_5638_), .B(_5613_), .Y(_5639_) );
NOR2X1 NOR2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_5638_), .B(_5613_), .Y(_5640_) );
INVX2 INVX2_194 ( .gnd(gnd), .vdd(vdd), .A(_5640_), .Y(_5641_) );
NAND3X1 NAND3X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_4850_), .B(_5639_), .C(_5641_), .Y(_5642_) );
INVX1 INVX1_750 ( .gnd(gnd), .vdd(vdd), .A(_5639_), .Y(_5643_) );
OAI21X1 OAI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(_5643_), .B(_5640_), .C(_4851_), .Y(_5644_) );
NAND3X1 NAND3X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_4854_), .B(_5644_), .C(_5642_), .Y(_5645_) );
NAND2X1 NAND2X1_754 ( .gnd(gnd), .vdd(vdd), .A(_5644_), .B(_5642_), .Y(_5646_) );
OAI21X1 OAI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(_4778_), .B(_4852_), .C(_5646_), .Y(_5647_) );
NAND2X1 NAND2X1_755 ( .gnd(gnd), .vdd(vdd), .A(_5645_), .B(_5647_), .Y(_5648_) );
INVX1 INVX1_751 ( .gnd(gnd), .vdd(vdd), .A(_5648_), .Y(_5649_) );
OAI21X1 OAI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(_5632_), .B(_5637_), .C(_5649_), .Y(_5650_) );
NAND3X1 NAND3X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_5634_), .B(_5635_), .C(_5636_), .Y(_5651_) );
AOI21X1 AOI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(_5630_), .B(_5629_), .C(_5136_), .Y(_5652_) );
AOI21X1 AOI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_5622_), .B(_5627_), .C(_5130_), .Y(_5653_) );
OAI21X1 OAI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(_5652_), .B(_5653_), .C(_5263_), .Y(_5654_) );
NAND3X1 NAND3X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_5648_), .B(_5651_), .C(_5654_), .Y(_5655_) );
NAND3X1 NAND3X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_5261_), .B(_5655_), .C(_5650_), .Y(_5656_) );
NAND2X1 NAND2X1_756 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_182_), .B(_5656_), .Y(_5657_) );
INVX2 INVX2_195 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_182_), .Y(_5658_) );
NAND3X1 NAND3X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_5649_), .B(_5651_), .C(_5654_), .Y(_5659_) );
OAI21X1 OAI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(_5632_), .B(_5637_), .C(_5648_), .Y(_5660_) );
AOI21X1 AOI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_5659_), .B(_5660_), .C(_7889_), .Y(_5661_) );
NAND2X1 NAND2X1_757 ( .gnd(gnd), .vdd(vdd), .A(_5658_), .B(_5661_), .Y(_5662_) );
NAND3X1 NAND3X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_5147_), .B(_5657_), .C(_5662_), .Y(_5663_) );
NAND2X1 NAND2X1_758 ( .gnd(gnd), .vdd(vdd), .A(_5659_), .B(_5660_), .Y(_5664_) );
NAND3X1 NAND3X1_1262 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_182_), .B(_5261_), .C(_5664_), .Y(_5665_) );
NAND2X1 NAND2X1_759 ( .gnd(gnd), .vdd(vdd), .A(_5658_), .B(_5656_), .Y(_5666_) );
NAND3X1 NAND3X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_5154_), .B(_5665_), .C(_5666_), .Y(_5667_) );
NAND3X1 NAND3X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_5667_), .B(_5260_), .C(_5663_), .Y(_5668_) );
AOI21X1 AOI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(_5147_), .B(_5152_), .C(_4657_), .Y(_5669_) );
AOI21X1 AOI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(_5160_), .B(_5158_), .C(_5669_), .Y(_5670_) );
AOI21X1 AOI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_5665_), .B(_5666_), .C(_5154_), .Y(_5671_) );
AOI21X1 AOI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_5657_), .B(_5662_), .C(_5147_), .Y(_5672_) );
OAI21X1 OAI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_5672_), .B(_5671_), .C(_5670_), .Y(_5673_) );
INVX1 INVX1_752 ( .gnd(gnd), .vdd(vdd), .A(_4863_), .Y(_5674_) );
INVX1 INVX1_753 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_170_), .Y(_5675_) );
NAND2X1 NAND2X1_760 ( .gnd(gnd), .vdd(vdd), .A(_5675_), .B(_5648_), .Y(_5676_) );
INVX1 INVX1_754 ( .gnd(gnd), .vdd(vdd), .A(_5676_), .Y(_5677_) );
NOR2X1 NOR2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_5675_), .B(_5648_), .Y(_5678_) );
NOR2X1 NOR2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_5678_), .B(_5677_), .Y(_5679_) );
AND2X2 AND2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_5679_), .B(_4860_), .Y(_5680_) );
OAI21X1 OAI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_5677_), .B(_5678_), .C(_4859_), .Y(_5681_) );
INVX1 INVX1_755 ( .gnd(gnd), .vdd(vdd), .A(_5681_), .Y(_5682_) );
NOR2X1 NOR2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_5682_), .B(_5680_), .Y(_5683_) );
NAND2X1 NAND2X1_761 ( .gnd(gnd), .vdd(vdd), .A(_5674_), .B(_5683_), .Y(_5684_) );
OAI21X1 OAI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(_5680_), .B(_5682_), .C(_4863_), .Y(_5685_) );
NAND2X1 NAND2X1_762 ( .gnd(gnd), .vdd(vdd), .A(_5685_), .B(_5684_), .Y(_5686_) );
NAND3X1 NAND3X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_5668_), .B(_5686_), .C(_5673_), .Y(_5687_) );
NAND3X1 NAND3X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_5154_), .B(_5657_), .C(_5662_), .Y(_5688_) );
NAND3X1 NAND3X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_5147_), .B(_5665_), .C(_5666_), .Y(_5689_) );
AOI21X1 AOI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(_5689_), .B(_5688_), .C(_5670_), .Y(_5690_) );
AOI21X1 AOI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_5667_), .B(_5663_), .C(_5260_), .Y(_5691_) );
INVX1 INVX1_756 ( .gnd(gnd), .vdd(vdd), .A(_5686_), .Y(_5692_) );
OAI21X1 OAI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(_5690_), .B(_5691_), .C(_5692_), .Y(_5693_) );
NAND3X1 NAND3X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_5258_), .B(_5687_), .C(_5693_), .Y(_5694_) );
NAND2X1 NAND2X1_763 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_198_), .B(_5694_), .Y(_5695_) );
INVX2 INVX2_196 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_198_), .Y(_5696_) );
AOI21X1 AOI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(_5668_), .B(_5673_), .C(_5686_), .Y(_5697_) );
NOR2X1 NOR2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_5257_), .B(_5697_), .Y(_5698_) );
NAND3X1 NAND3X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_5696_), .B(_5687_), .C(_5698_), .Y(_5699_) );
NAND3X1 NAND3X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_5173_), .B(_5695_), .C(_5699_), .Y(_5700_) );
NAND3X1 NAND3X1_1271 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_198_), .B(_5687_), .C(_5698_), .Y(_5701_) );
NAND2X1 NAND2X1_764 ( .gnd(gnd), .vdd(vdd), .A(_5696_), .B(_5694_), .Y(_5702_) );
NAND3X1 NAND3X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_5167_), .B(_5702_), .C(_5701_), .Y(_5703_) );
AOI21X1 AOI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(_5700_), .B(_5703_), .C(_5256_), .Y(_5704_) );
NOR3X1 NOR3X1_152 ( .gnd(gnd), .vdd(vdd), .A(_5174_), .B(_4906_), .C(_5173_), .Y(_5705_) );
OAI21X1 OAI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_5705_), .B(_4905_), .C(_5178_), .Y(_5706_) );
NAND3X1 NAND3X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_5167_), .B(_5695_), .C(_5699_), .Y(_5707_) );
NAND3X1 NAND3X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_5173_), .B(_5702_), .C(_5701_), .Y(_5708_) );
AOI21X1 AOI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_5707_), .B(_5708_), .C(_5706_), .Y(_5709_) );
INVX1 INVX1_757 ( .gnd(gnd), .vdd(vdd), .A(_4871_), .Y(_5710_) );
INVX1 INVX1_758 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_186_), .Y(_5711_) );
NAND2X1 NAND2X1_765 ( .gnd(gnd), .vdd(vdd), .A(_5711_), .B(_5686_), .Y(_5712_) );
NOR2X1 NOR2X1_442 ( .gnd(gnd), .vdd(vdd), .A(_5711_), .B(_5686_), .Y(_5713_) );
INVX1 INVX1_759 ( .gnd(gnd), .vdd(vdd), .A(_5713_), .Y(_5714_) );
NAND3X1 NAND3X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_4868_), .B(_5712_), .C(_5714_), .Y(_5715_) );
INVX1 INVX1_760 ( .gnd(gnd), .vdd(vdd), .A(_5712_), .Y(_5716_) );
OAI21X1 OAI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_5716_), .B(_5713_), .C(_4867_), .Y(_5717_) );
NAND3X1 NAND3X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_5710_), .B(_5717_), .C(_5715_), .Y(_5718_) );
INVX1 INVX1_761 ( .gnd(gnd), .vdd(vdd), .A(_5715_), .Y(_5719_) );
INVX1 INVX1_762 ( .gnd(gnd), .vdd(vdd), .A(_5717_), .Y(_5720_) );
OAI21X1 OAI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_5719_), .B(_5720_), .C(_4871_), .Y(_5721_) );
NAND2X1 NAND2X1_766 ( .gnd(gnd), .vdd(vdd), .A(_5718_), .B(_5721_), .Y(_5722_) );
INVX1 INVX1_763 ( .gnd(gnd), .vdd(vdd), .A(_5722_), .Y(_5723_) );
OAI21X1 OAI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5709_), .C(_5723_), .Y(_5724_) );
NAND3X1 NAND3X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_5707_), .B(_5708_), .C(_5706_), .Y(_5725_) );
AOI21X1 AOI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(_5702_), .B(_5701_), .C(_5173_), .Y(_5726_) );
AOI21X1 AOI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_5695_), .B(_5699_), .C(_5167_), .Y(_5727_) );
OAI21X1 OAI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(_5726_), .B(_5727_), .C(_5256_), .Y(_5728_) );
NAND3X1 NAND3X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_5725_), .B(_5722_), .C(_5728_), .Y(_5729_) );
NAND3X1 NAND3X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_5254_), .B(_5729_), .C(_5724_), .Y(_5730_) );
NAND2X1 NAND2X1_767 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_214_), .B(_5730_), .Y(_5731_) );
INVX2 INVX2_197 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_214_), .Y(_5732_) );
OAI21X1 OAI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5709_), .C(_5722_), .Y(_5733_) );
NAND3X1 NAND3X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_5725_), .B(_5723_), .C(_5728_), .Y(_5734_) );
AOI21X1 AOI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(_5734_), .B(_5733_), .C(_7907_), .Y(_5735_) );
NAND2X1 NAND2X1_768 ( .gnd(gnd), .vdd(vdd), .A(_5732_), .B(_5735_), .Y(_5736_) );
NAND3X1 NAND3X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_5192_), .B(_5731_), .C(_5736_), .Y(_5737_) );
NAND2X1 NAND2X1_769 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_214_), .B(_5735_), .Y(_5738_) );
NAND2X1 NAND2X1_770 ( .gnd(gnd), .vdd(vdd), .A(_5732_), .B(_5730_), .Y(_5739_) );
NAND3X1 NAND3X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_5186_), .B(_5739_), .C(_5738_), .Y(_5740_) );
AOI21X1 AOI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_5737_), .B(_5740_), .C(_5253_), .Y(_5741_) );
NOR3X1 NOR3X1_153 ( .gnd(gnd), .vdd(vdd), .A(_5193_), .B(_4903_), .C(_5192_), .Y(_5742_) );
OAI21X1 OAI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_5742_), .B(_4902_), .C(_5197_), .Y(_5743_) );
NAND3X1 NAND3X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_5186_), .B(_5731_), .C(_5736_), .Y(_5744_) );
NAND3X1 NAND3X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_5192_), .B(_5739_), .C(_5738_), .Y(_5745_) );
AOI21X1 AOI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_5744_), .B(_5745_), .C(_5743_), .Y(_5746_) );
INVX1 INVX1_764 ( .gnd(gnd), .vdd(vdd), .A(_4879_), .Y(_5747_) );
INVX1 INVX1_765 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_202_), .Y(_5748_) );
NAND2X1 NAND2X1_771 ( .gnd(gnd), .vdd(vdd), .A(_5748_), .B(_5722_), .Y(_5749_) );
NOR2X1 NOR2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_5748_), .B(_5722_), .Y(_5750_) );
INVX2 INVX2_198 ( .gnd(gnd), .vdd(vdd), .A(_5750_), .Y(_5751_) );
NAND3X1 NAND3X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_4876_), .B(_5749_), .C(_5751_), .Y(_5752_) );
INVX1 INVX1_766 ( .gnd(gnd), .vdd(vdd), .A(_5749_), .Y(_5753_) );
OAI21X1 OAI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_5753_), .B(_5750_), .C(_4875_), .Y(_5754_) );
NAND3X1 NAND3X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_5747_), .B(_5754_), .C(_5752_), .Y(_5755_) );
INVX1 INVX1_767 ( .gnd(gnd), .vdd(vdd), .A(_5752_), .Y(_5756_) );
INVX1 INVX1_768 ( .gnd(gnd), .vdd(vdd), .A(_5754_), .Y(_5757_) );
OAI21X1 OAI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_5756_), .B(_5757_), .C(_4879_), .Y(_5758_) );
NAND2X1 NAND2X1_772 ( .gnd(gnd), .vdd(vdd), .A(_5755_), .B(_5758_), .Y(_5759_) );
INVX2 INVX2_199 ( .gnd(gnd), .vdd(vdd), .A(_5759_), .Y(_5760_) );
OAI21X1 OAI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_5746_), .B(_5741_), .C(_5760_), .Y(_5761_) );
NAND3X1 NAND3X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_5744_), .B(_5745_), .C(_5743_), .Y(_5762_) );
AOI21X1 AOI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(_5739_), .B(_5738_), .C(_5192_), .Y(_5763_) );
AOI21X1 AOI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_5731_), .B(_5736_), .C(_5186_), .Y(_5764_) );
OAI21X1 OAI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_5763_), .B(_5764_), .C(_5253_), .Y(_5765_) );
NAND3X1 NAND3X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_5759_), .B(_5765_), .C(_5762_), .Y(_5766_) );
NAND3X1 NAND3X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_5251_), .B(_5766_), .C(_5761_), .Y(_5767_) );
NAND2X1 NAND2X1_773 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_230_), .B(_5767_), .Y(_5768_) );
INVX2 INVX2_200 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_230_), .Y(_5769_) );
OAI21X1 OAI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_5746_), .B(_5741_), .C(_5759_), .Y(_5770_) );
NAND3X1 NAND3X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_5760_), .B(_5765_), .C(_5762_), .Y(_5771_) );
AOI21X1 AOI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_5771_), .B(_5770_), .C(_5250_), .Y(_5772_) );
NAND2X1 NAND2X1_774 ( .gnd(gnd), .vdd(vdd), .A(_5769_), .B(_5772_), .Y(_5773_) );
NAND3X1 NAND3X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_5211_), .B(_5768_), .C(_5773_), .Y(_5774_) );
NAND2X1 NAND2X1_775 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_230_), .B(_5772_), .Y(_5775_) );
NAND2X1 NAND2X1_776 ( .gnd(gnd), .vdd(vdd), .A(_5769_), .B(_5767_), .Y(_5776_) );
NAND3X1 NAND3X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_5205_), .B(_5776_), .C(_5775_), .Y(_5777_) );
AOI21X1 AOI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(_5774_), .B(_5777_), .C(_5247_), .Y(_5778_) );
NOR3X1 NOR3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_5212_), .B(_4900_), .C(_5211_), .Y(_5779_) );
OAI21X1 OAI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(_5779_), .B(_4899_), .C(_5216_), .Y(_5780_) );
NAND3X1 NAND3X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_5205_), .B(_5768_), .C(_5773_), .Y(_5781_) );
NAND3X1 NAND3X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_5211_), .B(_5776_), .C(_5775_), .Y(_5782_) );
AOI21X1 AOI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(_5781_), .B(_5782_), .C(_5780_), .Y(_5783_) );
INVX1 INVX1_769 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .Y(_5784_) );
INVX1 INVX1_770 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_218_), .Y(_5785_) );
NAND2X1 NAND2X1_777 ( .gnd(gnd), .vdd(vdd), .A(_5785_), .B(_5759_), .Y(_5786_) );
NOR2X1 NOR2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_5785_), .B(_5759_), .Y(_5787_) );
INVX2 INVX2_201 ( .gnd(gnd), .vdd(vdd), .A(_5787_), .Y(_5788_) );
NAND2X1 NAND2X1_778 ( .gnd(gnd), .vdd(vdd), .A(_5786_), .B(_5788_), .Y(_5789_) );
OR2X2 OR2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_5789_), .B(_4883_), .Y(_5790_) );
AOI21X1 AOI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(_5786_), .B(_5788_), .C(_4884_), .Y(_5791_) );
INVX1 INVX1_771 ( .gnd(gnd), .vdd(vdd), .A(_5791_), .Y(_5792_) );
NAND3X1 NAND3X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_5784_), .B(_5792_), .C(_5790_), .Y(_5793_) );
NOR2X1 NOR2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_4883_), .B(_5789_), .Y(_5794_) );
OAI21X1 OAI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_5794_), .B(_5791_), .C(_4887_), .Y(_5795_) );
NAND2X1 NAND2X1_779 ( .gnd(gnd), .vdd(vdd), .A(_5795_), .B(_5793_), .Y(_5796_) );
INVX2 INVX2_202 ( .gnd(gnd), .vdd(vdd), .A(_5796_), .Y(_5797_) );
OAI21X1 OAI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_5783_), .B(_5778_), .C(_5797_), .Y(_5798_) );
NAND3X1 NAND3X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_5781_), .B(_5782_), .C(_5780_), .Y(_5799_) );
AOI21X1 AOI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_5776_), .B(_5775_), .C(_5211_), .Y(_5800_) );
AOI21X1 AOI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_5768_), .B(_5773_), .C(_5205_), .Y(_5801_) );
OAI21X1 OAI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_5800_), .B(_5801_), .C(_5247_), .Y(_5802_) );
NAND3X1 NAND3X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_5802_), .B(_5796_), .C(_5799_), .Y(_5803_) );
NAND3X1 NAND3X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_8157_), .B(_5803_), .C(_5798_), .Y(_5804_) );
NAND2X1 NAND2X1_780 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_246_), .B(_5804_), .Y(_5805_) );
INVX1 INVX1_772 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_246_), .Y(_5806_) );
NAND3X1 NAND3X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_5802_), .B(_5797_), .C(_5799_), .Y(_5807_) );
OAI21X1 OAI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(_5783_), .B(_5778_), .C(_5796_), .Y(_5808_) );
AOI21X1 AOI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(_5807_), .B(_5808_), .C(_7929_), .Y(_5809_) );
NAND2X1 NAND2X1_781 ( .gnd(gnd), .vdd(vdd), .A(_5806_), .B(_5809_), .Y(_5810_) );
NAND3X1 NAND3X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_5230_), .B(_5805_), .C(_5810_), .Y(_5811_) );
NAND2X1 NAND2X1_782 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_246_), .B(_5809_), .Y(_5812_) );
NAND2X1 NAND2X1_783 ( .gnd(gnd), .vdd(vdd), .A(_5806_), .B(_5804_), .Y(_5813_) );
NAND3X1 NAND3X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_5222_), .B(_5813_), .C(_5812_), .Y(_5814_) );
AOI21X1 AOI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(_5811_), .B(_5814_), .C(_5245_), .Y(_5815_) );
OAI21X1 OAI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_5235_), .B(_5234_), .C(_5232_), .Y(_5816_) );
NAND3X1 NAND3X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_5222_), .B(_5805_), .C(_5810_), .Y(_5817_) );
NAND3X1 NAND3X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_5230_), .B(_5813_), .C(_5812_), .Y(_5818_) );
AOI21X1 AOI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(_5817_), .B(_5818_), .C(_5816_), .Y(_5819_) );
INVX1 INVX1_773 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_5820_) );
NOR2X1 NOR2X1_446 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_234_), .B(_5797_), .Y(_5821_) );
INVX1 INVX1_774 ( .gnd(gnd), .vdd(vdd), .A(_5821_), .Y(_5822_) );
NAND2X1 NAND2X1_784 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_234_), .B(_5797_), .Y(_5823_) );
NAND3X1 NAND3X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_4892_), .B(_5823_), .C(_5822_), .Y(_5824_) );
INVX2 INVX2_203 ( .gnd(gnd), .vdd(vdd), .A(_5823_), .Y(_5825_) );
OAI21X1 OAI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(_5825_), .B(_5821_), .C(_4891_), .Y(_5826_) );
NAND3X1 NAND3X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_5820_), .B(_5826_), .C(_5824_), .Y(_5827_) );
NOR3X1 NOR3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_4891_), .B(_5821_), .C(_5825_), .Y(_5828_) );
AOI21X1 AOI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(_5823_), .B(_5822_), .C(_4892_), .Y(_5829_) );
OAI21X1 OAI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(_5829_), .B(_5828_), .C(_4895_), .Y(_5830_) );
NAND2X1 NAND2X1_785 ( .gnd(gnd), .vdd(vdd), .A(_5827_), .B(_5830_), .Y(_5831_) );
INVX2 INVX2_204 ( .gnd(gnd), .vdd(vdd), .A(_5831_), .Y(_5832_) );
OAI21X1 OAI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_5819_), .B(_5815_), .C(_5832_), .Y(_5833_) );
NAND3X1 NAND3X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_5817_), .B(_5818_), .C(_5816_), .Y(_5834_) );
NAND3X1 NAND3X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_5811_), .B(_5814_), .C(_5245_), .Y(_5835_) );
NAND3X1 NAND3X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_5835_), .B(_5831_), .C(_5834_), .Y(_5836_) );
NAND2X1 NAND2X1_786 ( .gnd(gnd), .vdd(vdd), .A(_5836_), .B(_5833_), .Y(_5837_) );
XOR2X1 XOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_5837_), .B(_5244_), .Y(module_1_H_6_) );
OAI21X1 OAI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(_5819_), .B(_5815_), .C(_5831_), .Y(_5838_) );
NAND3X1 NAND3X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_5835_), .B(_5832_), .C(_5834_), .Y(_5839_) );
NAND3X1 NAND3X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_5839_), .B(_5838_), .C(_5244_), .Y(_5840_) );
AOI21X1 AOI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_5813_), .B(_5812_), .C(_5230_), .Y(_5841_) );
AOI21X1 AOI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_5818_), .B(_5816_), .C(_5841_), .Y(_5842_) );
AOI21X1 AOI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_5820_), .B(_5826_), .C(_5828_), .Y(_5843_) );
OAI21X1 OAI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_5791_), .C(_5790_), .Y(_5844_) );
AOI21X1 AOI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_5747_), .B(_5754_), .C(_5756_), .Y(_5845_) );
INVX1 INVX1_775 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_203_), .Y(_5846_) );
OAI21X1 OAI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_5720_), .B(_4871_), .C(_5715_), .Y(_5847_) );
INVX1 INVX1_776 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_187_), .Y(_5848_) );
AOI21X1 AOI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_5674_), .B(_5681_), .C(_5680_), .Y(_5849_) );
INVX1 INVX1_777 ( .gnd(gnd), .vdd(vdd), .A(_5849_), .Y(_5850_) );
INVX1 INVX1_778 ( .gnd(gnd), .vdd(vdd), .A(_5678_), .Y(_5851_) );
INVX1 INVX1_779 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_171_), .Y(_5852_) );
OAI21X1 OAI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_5646_), .B(_4855_), .C(_5642_), .Y(_5853_) );
INVX1 INVX1_780 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_155_), .Y(_5854_) );
AOI21X1 AOI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_4846_), .B(_5609_), .C(_5607_), .Y(_5855_) );
INVX1 INVX1_781 ( .gnd(gnd), .vdd(vdd), .A(_5573_), .Y(_5856_) );
OAI21X1 OAI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_5856_), .B(_4839_), .C(_5570_), .Y(_5857_) );
OAI21X1 OAI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_4832_), .B(_5532_), .C(_5535_), .Y(_5858_) );
INVX1 INVX1_782 ( .gnd(gnd), .vdd(vdd), .A(_5528_), .Y(_5859_) );
OAI21X1 OAI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_4826_), .B(_5492_), .C(_5495_), .Y(_5860_) );
AOI21X1 AOI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_5453_), .B(_5455_), .C(_5448_), .Y(_5861_) );
INVX1 INVX1_783 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf2_), .Y(_5862_) );
NOR2X1 NOR2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_4788_), .B(_4809_), .Y(_5863_) );
AOI21X1 AOI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_5863_), .B(_5412_), .C(_5415_), .Y(_5864_) );
INVX1 INVX1_784 ( .gnd(gnd), .vdd(vdd), .A(_5376_), .Y(_5865_) );
AOI21X1 AOI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(_5369_), .B(_5865_), .C(_5375_), .Y(_5866_) );
INVX1 INVX1_785 ( .gnd(gnd), .vdd(vdd), .A(_5373_), .Y(_5867_) );
INVX1 INVX1_786 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .Y(_5868_) );
OAI21X1 OAI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_5343_), .B(_5340_), .C(_5336_), .Y(_5869_) );
NOR2X1 NOR2X1_448 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_27_), .B(module_1_W_11_), .Y(_5870_) );
INVX1 INVX1_787 ( .gnd(gnd), .vdd(vdd), .A(_5870_), .Y(_5871_) );
NAND2X1 NAND2X1_787 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_27_), .B(module_1_W_11_), .Y(_5872_) );
NAND2X1 NAND2X1_788 ( .gnd(gnd), .vdd(vdd), .A(_5872_), .B(_5871_), .Y(_5873_) );
NAND3X1 NAND3X1_1311 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_26_), .B(module_1_W_10_), .C(_5873_), .Y(_5874_) );
NAND3X1 NAND3X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_5332_), .B(_5872_), .C(_5871_), .Y(_5875_) );
NAND2X1 NAND2X1_789 ( .gnd(gnd), .vdd(vdd), .A(_5875_), .B(_5874_), .Y(_5876_) );
XOR2X1 XOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_5869_), .B(_5876_), .Y(_5877_) );
NAND2X1 NAND2X1_790 ( .gnd(gnd), .vdd(vdd), .A(_5868_), .B(_5877_), .Y(_5878_) );
XNOR2X1 XNOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_5869_), .B(_5876_), .Y(_5879_) );
NAND2X1 NAND2X1_791 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .B(_5879_), .Y(_5880_) );
NAND2X1 NAND2X1_792 ( .gnd(gnd), .vdd(vdd), .A(_5880_), .B(_5878_), .Y(_5881_) );
NAND2X1 NAND2X1_793 ( .gnd(gnd), .vdd(vdd), .A(_5867_), .B(_5881_), .Y(_5882_) );
NAND3X1 NAND3X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_5373_), .B(_5880_), .C(_5878_), .Y(_5883_) );
NAND2X1 NAND2X1_794 ( .gnd(gnd), .vdd(vdd), .A(_5883_), .B(_5882_), .Y(_5884_) );
XNOR2X1 XNOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_5884_), .B(_5866_), .Y(_5885_) );
NAND2X1 NAND2X1_795 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf2_), .B(_5885_), .Y(_5886_) );
INVX1 INVX1_788 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf1_), .Y(_5887_) );
OR2X2 OR2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_5374_), .B(_5370_), .Y(_5888_) );
OAI21X1 OAI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_4804_), .B(_5376_), .C(_5888_), .Y(_5889_) );
XNOR2X1 XNOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_5884_), .B(_5889_), .Y(_5890_) );
NAND2X1 NAND2X1_796 ( .gnd(gnd), .vdd(vdd), .A(_5887_), .B(_5890_), .Y(_5891_) );
NAND2X1 NAND2X1_797 ( .gnd(gnd), .vdd(vdd), .A(_5886_), .B(_5891_), .Y(_5892_) );
NOR2X1 NOR2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_5407_), .B(_5892_), .Y(_5893_) );
AOI21X1 AOI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_5886_), .B(_5891_), .C(_5411_), .Y(_5894_) );
OAI21X1 OAI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_5893_), .B(_5894_), .C(_5864_), .Y(_5895_) );
OAI21X1 OAI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(_5416_), .B(_4810_), .C(_5408_), .Y(_5896_) );
OR2X2 OR2X2_129 ( .gnd(gnd), .vdd(vdd), .A(_5892_), .B(_5407_), .Y(_5897_) );
INVX1 INVX1_789 ( .gnd(gnd), .vdd(vdd), .A(_5894_), .Y(_5898_) );
NAND3X1 NAND3X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_5898_), .B(_5896_), .C(_5897_), .Y(_5899_) );
NAND2X1 NAND2X1_798 ( .gnd(gnd), .vdd(vdd), .A(_5895_), .B(_5899_), .Y(_5900_) );
NAND2X1 NAND2X1_799 ( .gnd(gnd), .vdd(vdd), .A(_5862_), .B(_5900_), .Y(_5901_) );
AND2X2 AND2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_5899_), .B(_5895_), .Y(_5902_) );
NAND2X1 NAND2X1_800 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf1_), .B(_5902_), .Y(_5903_) );
AOI21X1 AOI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_5901_), .B(_5903_), .C(_5450_), .Y(_5904_) );
NAND3X1 NAND3X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_5450_), .B(_5901_), .C(_5903_), .Y(_5905_) );
INVX2 INVX2_205 ( .gnd(gnd), .vdd(vdd), .A(_5905_), .Y(_5906_) );
OAI21X1 OAI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_5906_), .B(_5904_), .C(_5861_), .Y(_5907_) );
INVX2 INVX2_206 ( .gnd(gnd), .vdd(vdd), .A(_5907_), .Y(_5908_) );
NOR2X1 NOR2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_5904_), .B(_5906_), .Y(_5909_) );
OAI21X1 OAI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(_5448_), .B(_5452_), .C(_5909_), .Y(_5910_) );
INVX2 INVX2_207 ( .gnd(gnd), .vdd(vdd), .A(_5910_), .Y(_5911_) );
OAI21X1 OAI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(_5911_), .B(_5908_), .C(bloque_datos_59_bF_buf3_), .Y(_5912_) );
INVX1 INVX1_790 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf2_), .Y(_5913_) );
NAND3X1 NAND3X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_5913_), .B(_5907_), .C(_5910_), .Y(_5914_) );
NAND3X1 NAND3X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_5488_), .B(_5914_), .C(_5912_), .Y(_5915_) );
OAI21X1 OAI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_5911_), .B(_5908_), .C(_5913_), .Y(_5916_) );
NAND3X1 NAND3X1_1318 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf1_), .B(_5907_), .C(_5910_), .Y(_5917_) );
NAND3X1 NAND3X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_5491_), .B(_5917_), .C(_5916_), .Y(_5918_) );
AOI21X1 AOI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_5915_), .B(_5918_), .C(_5860_), .Y(_5919_) );
NAND3X1 NAND3X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_5860_), .B(_5915_), .C(_5918_), .Y(_5920_) );
INVX2 INVX2_208 ( .gnd(gnd), .vdd(vdd), .A(_5920_), .Y(_5921_) );
OAI21X1 OAI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(_5921_), .B(_5919_), .C(bloque_datos_75_bF_buf2_), .Y(_5922_) );
INVX1 INVX1_791 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf1_), .Y(_5923_) );
INVX1 INVX1_792 ( .gnd(gnd), .vdd(vdd), .A(_5919_), .Y(_5924_) );
NAND3X1 NAND3X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_5923_), .B(_5920_), .C(_5924_), .Y(_5925_) );
NAND3X1 NAND3X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_5859_), .B(_5925_), .C(_5922_), .Y(_5926_) );
OAI21X1 OAI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_5921_), .B(_5919_), .C(_5923_), .Y(_5927_) );
NAND3X1 NAND3X1_1323 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf0_), .B(_5920_), .C(_5924_), .Y(_5928_) );
NAND3X1 NAND3X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_5528_), .B(_5928_), .C(_5927_), .Y(_5929_) );
AOI21X1 AOI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(_5926_), .B(_5929_), .C(_5858_), .Y(_5930_) );
NAND3X1 NAND3X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_5858_), .B(_5926_), .C(_5929_), .Y(_5931_) );
INVX2 INVX2_209 ( .gnd(gnd), .vdd(vdd), .A(_5931_), .Y(_5932_) );
OAI21X1 OAI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(_5932_), .B(_5930_), .C(bloque_datos_91_bF_buf2_), .Y(_5933_) );
INVX1 INVX1_793 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf1_), .Y(_5934_) );
INVX1 INVX1_794 ( .gnd(gnd), .vdd(vdd), .A(_5930_), .Y(_5935_) );
NAND3X1 NAND3X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_5934_), .B(_5931_), .C(_5935_), .Y(_5936_) );
NAND3X1 NAND3X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_5572_), .B(_5936_), .C(_5933_), .Y(_5937_) );
OAI21X1 OAI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(_5932_), .B(_5930_), .C(_5934_), .Y(_5938_) );
NAND3X1 NAND3X1_1328 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf0_), .B(_5931_), .C(_5935_), .Y(_5939_) );
NAND3X1 NAND3X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_5569_), .B(_5939_), .C(_5938_), .Y(_5940_) );
NAND3X1 NAND3X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_5937_), .B(_5940_), .C(_5857_), .Y(_5941_) );
INVX1 INVX1_795 ( .gnd(gnd), .vdd(vdd), .A(_5941_), .Y(_5942_) );
AOI21X1 AOI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(_5937_), .B(_5940_), .C(_5857_), .Y(_5943_) );
NOR2X1 NOR2X1_451 ( .gnd(gnd), .vdd(vdd), .A(_5943_), .B(_5942_), .Y(_5944_) );
XNOR2X1 XNOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_5944_), .B(module_1_W_139_), .Y(_5945_) );
NOR2X1 NOR2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_5605_), .B(_5945_), .Y(_5946_) );
INVX1 INVX1_796 ( .gnd(gnd), .vdd(vdd), .A(_5946_), .Y(_5947_) );
OAI21X1 OAI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_5603_), .B(_5579_), .C(_5945_), .Y(_5948_) );
NAND2X1 NAND2X1_801 ( .gnd(gnd), .vdd(vdd), .A(_5948_), .B(_5947_), .Y(_5949_) );
OR2X2 OR2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_5949_), .B(_5855_), .Y(_5950_) );
INVX1 INVX1_797 ( .gnd(gnd), .vdd(vdd), .A(_5948_), .Y(_5951_) );
OAI21X1 OAI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_5951_), .B(_5946_), .C(_5855_), .Y(_5952_) );
NAND2X1 NAND2X1_802 ( .gnd(gnd), .vdd(vdd), .A(_5952_), .B(_5950_), .Y(_5953_) );
NAND2X1 NAND2X1_803 ( .gnd(gnd), .vdd(vdd), .A(_5854_), .B(_5953_), .Y(_5954_) );
INVX1 INVX1_798 ( .gnd(gnd), .vdd(vdd), .A(_5954_), .Y(_5955_) );
NOR2X1 NOR2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_5854_), .B(_5953_), .Y(_5956_) );
NOR3X1 NOR3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_5641_), .B(_5956_), .C(_5955_), .Y(_5957_) );
INVX2 INVX2_210 ( .gnd(gnd), .vdd(vdd), .A(_5956_), .Y(_5958_) );
AOI21X1 AOI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_5954_), .B(_5958_), .C(_5640_), .Y(_5959_) );
NOR2X1 NOR2X1_454 ( .gnd(gnd), .vdd(vdd), .A(_5957_), .B(_5959_), .Y(_5960_) );
AND2X2 AND2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_5960_), .B(_5853_), .Y(_5961_) );
AND2X2 AND2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_5645_), .B(_5642_), .Y(_5962_) );
OAI21X1 OAI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(_5959_), .B(_5957_), .C(_5962_), .Y(_5963_) );
INVX2 INVX2_211 ( .gnd(gnd), .vdd(vdd), .A(_5963_), .Y(_5964_) );
OAI21X1 OAI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(_5961_), .B(_5964_), .C(_5852_), .Y(_5965_) );
NOR2X1 NOR2X1_455 ( .gnd(gnd), .vdd(vdd), .A(_5964_), .B(_5961_), .Y(_5966_) );
NAND2X1 NAND2X1_804 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_171_), .B(_5966_), .Y(_5967_) );
NAND2X1 NAND2X1_805 ( .gnd(gnd), .vdd(vdd), .A(_5965_), .B(_5967_), .Y(_5968_) );
NOR2X1 NOR2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_5851_), .B(_5968_), .Y(_5969_) );
AOI21X1 AOI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(_5965_), .B(_5967_), .C(_5678_), .Y(_5970_) );
NOR2X1 NOR2X1_457 ( .gnd(gnd), .vdd(vdd), .A(_5970_), .B(_5969_), .Y(_5971_) );
AND2X2 AND2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_5971_), .B(_5850_), .Y(_5972_) );
OAI21X1 OAI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_5969_), .B(_5970_), .C(_5849_), .Y(_5973_) );
INVX2 INVX2_212 ( .gnd(gnd), .vdd(vdd), .A(_5973_), .Y(_5974_) );
OAI21X1 OAI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(_5972_), .B(_5974_), .C(_5848_), .Y(_5975_) );
NOR2X1 NOR2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_5974_), .B(_5972_), .Y(_5976_) );
NAND2X1 NAND2X1_806 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_187_), .B(_5976_), .Y(_5977_) );
NAND3X1 NAND3X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_5713_), .B(_5975_), .C(_5977_), .Y(_5978_) );
INVX2 INVX2_213 ( .gnd(gnd), .vdd(vdd), .A(_5978_), .Y(_5979_) );
AOI21X1 AOI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(_5975_), .B(_5977_), .C(_5713_), .Y(_5980_) );
NOR2X1 NOR2X1_459 ( .gnd(gnd), .vdd(vdd), .A(_5980_), .B(_5979_), .Y(_5981_) );
NAND2X1 NAND2X1_807 ( .gnd(gnd), .vdd(vdd), .A(_5847_), .B(_5981_), .Y(_5982_) );
AOI21X1 AOI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_5710_), .B(_5717_), .C(_5719_), .Y(_5983_) );
OAI21X1 OAI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_5979_), .B(_5980_), .C(_5983_), .Y(_5984_) );
NAND2X1 NAND2X1_808 ( .gnd(gnd), .vdd(vdd), .A(_5984_), .B(_5982_), .Y(_5985_) );
NAND2X1 NAND2X1_809 ( .gnd(gnd), .vdd(vdd), .A(_5846_), .B(_5985_), .Y(_5986_) );
NOR2X1 NOR2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_5846_), .B(_5985_), .Y(_5987_) );
INVX2 INVX2_214 ( .gnd(gnd), .vdd(vdd), .A(_5987_), .Y(_5988_) );
NAND3X1 NAND3X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_5750_), .B(_5986_), .C(_5988_), .Y(_5989_) );
INVX1 INVX1_799 ( .gnd(gnd), .vdd(vdd), .A(_5986_), .Y(_5990_) );
OAI21X1 OAI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(_5990_), .B(_5987_), .C(_5751_), .Y(_5991_) );
NAND2X1 NAND2X1_810 ( .gnd(gnd), .vdd(vdd), .A(_5991_), .B(_5989_), .Y(_5992_) );
NOR2X1 NOR2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_5845_), .B(_5992_), .Y(_5993_) );
OAI21X1 OAI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(_5757_), .B(_4879_), .C(_5752_), .Y(_5994_) );
AOI21X1 AOI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_5991_), .B(_5989_), .C(_5994_), .Y(_5995_) );
NOR2X1 NOR2X1_462 ( .gnd(gnd), .vdd(vdd), .A(_5995_), .B(_5993_), .Y(_5996_) );
NOR2X1 NOR2X1_463 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_219_), .B(_5996_), .Y(_5997_) );
AND2X2 AND2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_5996_), .B(module_1_W_219_), .Y(_5998_) );
NOR3X1 NOR3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_5997_), .B(_5788_), .C(_5998_), .Y(_5999_) );
OR2X2 OR2X2_131 ( .gnd(gnd), .vdd(vdd), .A(_5996_), .B(module_1_W_219_), .Y(_6000_) );
NAND2X1 NAND2X1_811 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_219_), .B(_5996_), .Y(_6001_) );
AOI21X1 AOI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_6001_), .B(_6000_), .C(_5787_), .Y(_6002_) );
NOR2X1 NOR2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_6002_), .B(_5999_), .Y(_6003_) );
AND2X2 AND2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_6003_), .B(_5844_), .Y(_6004_) );
NOR2X1 NOR2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_5844_), .B(_6003_), .Y(_6005_) );
NOR2X1 NOR2X1_466 ( .gnd(gnd), .vdd(vdd), .A(_6005_), .B(_6004_), .Y(_6006_) );
OR2X2 OR2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_6006_), .B(module_1_W_235_), .Y(_6007_) );
NAND2X1 NAND2X1_812 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_235_), .B(_6006_), .Y(_6008_) );
NAND3X1 NAND3X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_5825_), .B(_6008_), .C(_6007_), .Y(_6009_) );
INVX2 INVX2_215 ( .gnd(gnd), .vdd(vdd), .A(_6009_), .Y(_6010_) );
AOI21X1 AOI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(_6008_), .B(_6007_), .C(_5825_), .Y(_6011_) );
OAI21X1 OAI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(_6010_), .B(_6011_), .C(_5843_), .Y(_6012_) );
INVX1 INVX1_800 ( .gnd(gnd), .vdd(vdd), .A(_6012_), .Y(_6013_) );
OAI21X1 OAI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(_5829_), .B(_4895_), .C(_5824_), .Y(_6014_) );
NOR2X1 NOR2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_6011_), .B(_6010_), .Y(_6015_) );
AND2X2 AND2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_6015_), .B(_6014_), .Y(_6016_) );
NOR2X1 NOR2X1_468 ( .gnd(gnd), .vdd(vdd), .A(_6013_), .B(_6016_), .Y(_6017_) );
INVX2 INVX2_216 ( .gnd(gnd), .vdd(vdd), .A(_6017_), .Y(_6018_) );
INVX1 INVX1_801 ( .gnd(gnd), .vdd(vdd), .A(_6006_), .Y(_6019_) );
AOI21X1 AOI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(_5708_), .B(_5706_), .C(_5726_), .Y(_6020_) );
OAI21X1 OAI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(_5672_), .B(_5670_), .C(_5663_), .Y(_6021_) );
INVX1 INVX1_802 ( .gnd(gnd), .vdd(vdd), .A(_6021_), .Y(_6022_) );
OR2X2 OR2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_5972_), .B(_5974_), .Y(_6023_) );
OAI21X1 OAI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(_5626_), .B(_5623_), .C(module_1_W_167_), .Y(_6024_) );
INVX1 INVX1_803 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_167_), .Y(_6025_) );
NAND3X1 NAND3X1_1334 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_166_), .B(_6025_), .C(_5621_), .Y(_6026_) );
OR2X2 OR2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_5961_), .B(_5964_), .Y(_6027_) );
INVX1 INVX1_804 ( .gnd(gnd), .vdd(vdd), .A(_5550_), .Y(_6028_) );
AOI21X1 AOI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(_5271_), .B(_5518_), .C(_5521_), .Y(_6029_) );
INVX1 INVX1_805 ( .gnd(gnd), .vdd(vdd), .A(_6029_), .Y(_6030_) );
NOR2X1 NOR2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_5930_), .B(_5932_), .Y(_6031_) );
OAI21X1 OAI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(_5479_), .B(_5481_), .C(_5474_), .Y(_6032_) );
NOR2X1 NOR2X1_470 ( .gnd(gnd), .vdd(vdd), .A(_5919_), .B(_5921_), .Y(_6033_) );
OAI21X1 OAI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(_5437_), .B(_5439_), .C(_5432_), .Y(_6034_) );
NOR2X1 NOR2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_5908_), .B(_5911_), .Y(_6035_) );
INVX1 INVX1_806 ( .gnd(gnd), .vdd(vdd), .A(_6035_), .Y(_6036_) );
AOI21X1 AOI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(_5397_), .B(_5277_), .C(_5400_), .Y(_6037_) );
AOI21X1 AOI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_5362_), .B(_5279_), .C(_5365_), .Y(_6038_) );
AOI21X1 AOI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_5282_), .B(_5324_), .C(_5328_), .Y(_6039_) );
INVX1 INVX1_807 ( .gnd(gnd), .vdd(vdd), .A(_5299_), .Y(_6040_) );
NOR2X1 NOR2X1_472 ( .gnd(gnd), .vdd(vdd), .A(_6040_), .B(_5304_), .Y(_6041_) );
XNOR2X1 XNOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_7_), .B(module_1_W_23_), .Y(_6042_) );
XOR2X1 XOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_7980_), .B(_6042_), .Y(_6043_) );
XNOR2X1 XNOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_5290_), .B(module_1_W_11_), .Y(_6044_) );
XNOR2X1 XNOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_6044_), .B(_6043_), .Y(_6045_) );
XNOR2X1 XNOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_6045_), .B(_5294_), .Y(_6046_) );
NAND2X1 NAND2X1_813 ( .gnd(gnd), .vdd(vdd), .A(_7988_), .B(_7990_), .Y(_6047_) );
XNOR2X1 XNOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_6047_), .B(bloque_datos[7]), .Y(_6048_) );
NOR2X1 NOR2X1_473 ( .gnd(gnd), .vdd(vdd), .A(_6046_), .B(_6048_), .Y(_6049_) );
AND2X2 AND2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_6048_), .B(_6046_), .Y(_6050_) );
NOR2X1 NOR2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_6049_), .B(_6050_), .Y(_6051_) );
NOR2X1 NOR2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_6041_), .B(_6051_), .Y(_6052_) );
AND2X2 AND2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_6051_), .B(_6041_), .Y(_6053_) );
OAI21X1 OAI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(_6053_), .B(_6052_), .C(_5877_), .Y(_6054_) );
OR2X2 OR2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_6051_), .B(_6041_), .Y(_6055_) );
NAND2X1 NAND2X1_814 ( .gnd(gnd), .vdd(vdd), .A(_6041_), .B(_6051_), .Y(_6056_) );
NAND3X1 NAND3X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_5879_), .B(_6056_), .C(_6055_), .Y(_6057_) );
AND2X2 AND2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_6057_), .B(_6054_), .Y(_6058_) );
AOI21X1 AOI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_5319_), .B(_5318_), .C(_5317_), .Y(_6059_) );
OAI21X1 OAI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(_8007_), .B(_8002_), .C(bloque_datos_23_bF_buf3_), .Y(_6060_) );
NAND2X1 NAND2X1_815 ( .gnd(gnd), .vdd(vdd), .A(_8004_), .B(_8003_), .Y(_6061_) );
OR2X2 OR2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_6061_), .B(bloque_datos_23_bF_buf2_), .Y(_6062_) );
NAND3X1 NAND3X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_6060_), .B(_6059_), .C(_6062_), .Y(_6063_) );
INVX1 INVX1_808 ( .gnd(gnd), .vdd(vdd), .A(_6060_), .Y(_6064_) );
NOR2X1 NOR2X1_476 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf1_), .B(_6061_), .Y(_6065_) );
OAI21X1 OAI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(_6065_), .B(_6064_), .C(_5316_), .Y(_6066_) );
AOI21X1 AOI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_6063_), .B(_6066_), .C(_6058_), .Y(_6067_) );
NAND2X1 NAND2X1_816 ( .gnd(gnd), .vdd(vdd), .A(_6054_), .B(_6057_), .Y(_6068_) );
NAND2X1 NAND2X1_817 ( .gnd(gnd), .vdd(vdd), .A(_6066_), .B(_6063_), .Y(_6069_) );
NOR2X1 NOR2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_6068_), .B(_6069_), .Y(_6070_) );
OAI21X1 OAI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(_6070_), .B(_6067_), .C(_6039_), .Y(_6071_) );
INVX1 INVX1_809 ( .gnd(gnd), .vdd(vdd), .A(_6039_), .Y(_6072_) );
NOR3X1 NOR3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_6065_), .B(_6064_), .C(_5316_), .Y(_6073_) );
AOI21X1 AOI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_6060_), .B(_6062_), .C(_6059_), .Y(_6074_) );
OAI21X1 OAI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_6073_), .B(_6074_), .C(_6068_), .Y(_6075_) );
NAND3X1 NAND3X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_6063_), .B(_6066_), .C(_6058_), .Y(_6076_) );
NAND3X1 NAND3X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_6075_), .B(_6076_), .C(_6072_), .Y(_6077_) );
NAND3X1 NAND3X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_5885_), .B(_6077_), .C(_6071_), .Y(_6078_) );
OAI21X1 OAI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(_6070_), .B(_6067_), .C(_6072_), .Y(_6079_) );
NAND3X1 NAND3X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_6039_), .B(_6075_), .C(_6076_), .Y(_6080_) );
NAND3X1 NAND3X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_5890_), .B(_6080_), .C(_6079_), .Y(_6081_) );
NAND2X1 NAND2X1_818 ( .gnd(gnd), .vdd(vdd), .A(_6081_), .B(_6078_), .Y(_6082_) );
NAND2X1 NAND2X1_819 ( .gnd(gnd), .vdd(vdd), .A(_8021_), .B(_8020_), .Y(_6083_) );
XNOR2X1 XNOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_6083_), .B(bloque_datos[39]), .Y(_6084_) );
NOR2X1 NOR2X1_478 ( .gnd(gnd), .vdd(vdd), .A(_5354_), .B(_6084_), .Y(_6085_) );
AND2X2 AND2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_6084_), .B(_5354_), .Y(_6086_) );
OAI21X1 OAI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_6086_), .B(_6085_), .C(_6082_), .Y(_6087_) );
AND2X2 AND2X2_129 ( .gnd(gnd), .vdd(vdd), .A(_6078_), .B(_6081_), .Y(_6088_) );
OR2X2 OR2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_6084_), .B(_5354_), .Y(_6089_) );
NAND2X1 NAND2X1_820 ( .gnd(gnd), .vdd(vdd), .A(_5354_), .B(_6084_), .Y(_6090_) );
NAND3X1 NAND3X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_6089_), .B(_6090_), .C(_6088_), .Y(_6091_) );
NAND3X1 NAND3X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_6038_), .B(_6087_), .C(_6091_), .Y(_6092_) );
OAI21X1 OAI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(_5364_), .B(_5366_), .C(_5359_), .Y(_6093_) );
AOI21X1 AOI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_6089_), .B(_6090_), .C(_6088_), .Y(_6094_) );
NOR3X1 NOR3X1_159 ( .gnd(gnd), .vdd(vdd), .A(_6085_), .B(_6086_), .C(_6082_), .Y(_6095_) );
OAI21X1 OAI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(_6094_), .B(_6095_), .C(_6093_), .Y(_6096_) );
NAND3X1 NAND3X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_5900_), .B(_6092_), .C(_6096_), .Y(_6097_) );
NAND3X1 NAND3X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_6093_), .B(_6087_), .C(_6091_), .Y(_6098_) );
OAI21X1 OAI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(_6094_), .B(_6095_), .C(_6038_), .Y(_6099_) );
NAND3X1 NAND3X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_5902_), .B(_6098_), .C(_6099_), .Y(_6100_) );
AND2X2 AND2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_6097_), .B(_6100_), .Y(_6101_) );
XNOR2X1 XNOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_8030_), .B(bloque_datos[55]), .Y(_6102_) );
OR2X2 OR2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_6102_), .B(_5389_), .Y(_6103_) );
NAND2X1 NAND2X1_821 ( .gnd(gnd), .vdd(vdd), .A(_5389_), .B(_6102_), .Y(_6104_) );
AOI21X1 AOI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(_6104_), .B(_6103_), .C(_6101_), .Y(_6105_) );
NAND2X1 NAND2X1_822 ( .gnd(gnd), .vdd(vdd), .A(_6097_), .B(_6100_), .Y(_6106_) );
NOR2X1 NOR2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_5389_), .B(_6102_), .Y(_6107_) );
AND2X2 AND2X2_131 ( .gnd(gnd), .vdd(vdd), .A(_6102_), .B(_5389_), .Y(_6108_) );
NOR3X1 NOR3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_6108_), .B(_6107_), .C(_6106_), .Y(_6109_) );
OAI21X1 OAI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(_6105_), .B(_6109_), .C(_6037_), .Y(_6110_) );
OAI21X1 OAI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(_5399_), .B(_5401_), .C(_5394_), .Y(_6111_) );
OAI21X1 OAI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(_6108_), .B(_6107_), .C(_6106_), .Y(_6112_) );
NAND3X1 NAND3X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_6104_), .B(_6103_), .C(_6101_), .Y(_6113_) );
NAND3X1 NAND3X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_6112_), .B(_6111_), .C(_6113_), .Y(_6114_) );
NAND3X1 NAND3X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_6036_), .B(_6114_), .C(_6110_), .Y(_6115_) );
OAI21X1 OAI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(_6105_), .B(_6109_), .C(_6111_), .Y(_6116_) );
NAND3X1 NAND3X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_6037_), .B(_6112_), .C(_6113_), .Y(_6117_) );
NAND3X1 NAND3X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_6035_), .B(_6117_), .C(_6116_), .Y(_6118_) );
AND2X2 AND2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_6115_), .B(_6118_), .Y(_6119_) );
OAI21X1 OAI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_8036_), .B(_8042_), .C(bloque_datos_71_bF_buf3_), .Y(_6120_) );
INVX1 INVX1_810 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf2_), .Y(_6121_) );
OAI21X1 OAI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(_8038_), .B(_8041_), .C(_8037_), .Y(_6122_) );
NAND3X1 NAND3X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_7967_), .B(_8035_), .C(_8032_), .Y(_6123_) );
NAND3X1 NAND3X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_6121_), .B(_6122_), .C(_6123_), .Y(_6124_) );
NAND2X1 NAND2X1_823 ( .gnd(gnd), .vdd(vdd), .A(_6124_), .B(_6120_), .Y(_6125_) );
OR2X2 OR2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_6125_), .B(_5427_), .Y(_6126_) );
NAND2X1 NAND2X1_824 ( .gnd(gnd), .vdd(vdd), .A(_5427_), .B(_6125_), .Y(_6127_) );
AOI21X1 AOI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_6126_), .B(_6127_), .C(_6119_), .Y(_6128_) );
NAND2X1 NAND2X1_825 ( .gnd(gnd), .vdd(vdd), .A(_6115_), .B(_6118_), .Y(_6129_) );
NOR2X1 NOR2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_5427_), .B(_6125_), .Y(_6130_) );
AND2X2 AND2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_6125_), .B(_5427_), .Y(_6131_) );
NOR3X1 NOR3X1_161 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_6130_), .C(_6129_), .Y(_6132_) );
OAI21X1 OAI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_6128_), .B(_6132_), .C(_6034_), .Y(_6133_) );
AOI21X1 AOI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(_5435_), .B(_5275_), .C(_5438_), .Y(_6134_) );
OAI21X1 OAI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_6130_), .C(_6129_), .Y(_6135_) );
NAND3X1 NAND3X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_6126_), .B(_6127_), .C(_6119_), .Y(_6136_) );
NAND3X1 NAND3X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_6134_), .B(_6135_), .C(_6136_), .Y(_6137_) );
AOI21X1 AOI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(_6137_), .B(_6133_), .C(_6033_), .Y(_6138_) );
INVX1 INVX1_811 ( .gnd(gnd), .vdd(vdd), .A(_6033_), .Y(_6139_) );
OAI21X1 OAI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_6128_), .B(_6132_), .C(_6134_), .Y(_6140_) );
NAND3X1 NAND3X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_6135_), .B(_6034_), .C(_6136_), .Y(_6141_) );
AOI21X1 AOI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_6141_), .B(_6140_), .C(_6139_), .Y(_6142_) );
OR2X2 OR2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_6138_), .B(_6142_), .Y(_6143_) );
NAND3X1 NAND3X1_1357 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf2_), .B(_8052_), .C(_8056_), .Y(_6144_) );
INVX1 INVX1_812 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf1_), .Y(_6145_) );
OAI21X1 OAI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_8053_), .B(_8051_), .C(_6145_), .Y(_6146_) );
NAND2X1 NAND2X1_826 ( .gnd(gnd), .vdd(vdd), .A(_6144_), .B(_6146_), .Y(_6147_) );
OR2X2 OR2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_6147_), .B(_5469_), .Y(_6148_) );
NAND2X1 NAND2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_5469_), .B(_6147_), .Y(_6149_) );
NAND3X1 NAND3X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_6148_), .B(_6149_), .C(_6143_), .Y(_6150_) );
NOR2X1 NOR2X1_481 ( .gnd(gnd), .vdd(vdd), .A(_6138_), .B(_6142_), .Y(_6151_) );
NOR2X1 NOR2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_5469_), .B(_6147_), .Y(_6152_) );
AND2X2 AND2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_6147_), .B(_5469_), .Y(_6153_) );
OAI21X1 OAI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(_6153_), .B(_6152_), .C(_6151_), .Y(_6154_) );
NAND3X1 NAND3X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_6154_), .B(_6032_), .C(_6150_), .Y(_6155_) );
AOI21X1 AOI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_5477_), .B(_5273_), .C(_5480_), .Y(_6156_) );
NOR3X1 NOR3X1_162 ( .gnd(gnd), .vdd(vdd), .A(_6153_), .B(_6152_), .C(_6151_), .Y(_6157_) );
AOI21X1 AOI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(_6149_), .B(_6148_), .C(_6143_), .Y(_6158_) );
OAI21X1 OAI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(_6157_), .B(_6158_), .C(_6156_), .Y(_6159_) );
AOI21X1 AOI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(_6155_), .B(_6159_), .C(_6031_), .Y(_6160_) );
INVX1 INVX1_813 ( .gnd(gnd), .vdd(vdd), .A(_6031_), .Y(_6161_) );
NAND3X1 NAND3X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_6156_), .B(_6154_), .C(_6150_), .Y(_6162_) );
OAI21X1 OAI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(_6157_), .B(_6158_), .C(_6032_), .Y(_6163_) );
AOI21X1 AOI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(_6162_), .B(_6163_), .C(_6161_), .Y(_6164_) );
NOR2X1 NOR2X1_483 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .B(_6164_), .Y(_6165_) );
NAND3X1 NAND3X1_1361 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_135_), .B(_8064_), .C(_8067_), .Y(_6166_) );
INVX1 INVX1_814 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_135_), .Y(_6167_) );
OAI21X1 OAI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(_8065_), .B(_8063_), .C(_6167_), .Y(_6168_) );
NAND2X1 NAND2X1_828 ( .gnd(gnd), .vdd(vdd), .A(_6166_), .B(_6168_), .Y(_6169_) );
NOR2X1 NOR2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_6169_), .B(_5510_), .Y(_6170_) );
NAND2X1 NAND2X1_829 ( .gnd(gnd), .vdd(vdd), .A(_6169_), .B(_5510_), .Y(_6171_) );
INVX1 INVX1_815 ( .gnd(gnd), .vdd(vdd), .A(_6171_), .Y(_6172_) );
NOR3X1 NOR3X1_163 ( .gnd(gnd), .vdd(vdd), .A(_6172_), .B(_6170_), .C(_6165_), .Y(_6173_) );
OR2X2 OR2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .B(_6164_), .Y(_6174_) );
INVX1 INVX1_816 ( .gnd(gnd), .vdd(vdd), .A(_6170_), .Y(_6175_) );
AOI21X1 AOI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(_6171_), .B(_6175_), .C(_6174_), .Y(_6176_) );
OAI21X1 OAI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(_6173_), .B(_6176_), .C(_6030_), .Y(_6177_) );
NAND3X1 NAND3X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_6171_), .B(_6175_), .C(_6174_), .Y(_6178_) );
OAI21X1 OAI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(_6172_), .B(_6170_), .C(_6165_), .Y(_6179_) );
NAND3X1 NAND3X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_6029_), .B(_6179_), .C(_6178_), .Y(_6180_) );
AOI21X1 AOI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(_6180_), .B(_6177_), .C(_5944_), .Y(_6181_) );
INVX1 INVX1_817 ( .gnd(gnd), .vdd(vdd), .A(_5944_), .Y(_6182_) );
OAI21X1 OAI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_6173_), .B(_6176_), .C(_6029_), .Y(_6183_) );
NAND3X1 NAND3X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_6179_), .B(_6178_), .C(_6030_), .Y(_6184_) );
AOI21X1 AOI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(_6184_), .B(_6183_), .C(_6182_), .Y(_6185_) );
OAI21X1 OAI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(_6181_), .B(_6185_), .C(_6028_), .Y(_6186_) );
NAND3X1 NAND3X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_6182_), .B(_6184_), .C(_6183_), .Y(_6187_) );
NAND3X1 NAND3X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_5944_), .B(_6180_), .C(_6177_), .Y(_6188_) );
NAND3X1 NAND3X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_5550_), .B(_6187_), .C(_6188_), .Y(_6189_) );
NAND2X1 NAND2X1_830 ( .gnd(gnd), .vdd(vdd), .A(_6189_), .B(_6186_), .Y(_6190_) );
OAI21X1 OAI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(_5561_), .B(_5583_), .C(_6190_), .Y(_6191_) );
INVX1 INVX1_818 ( .gnd(gnd), .vdd(vdd), .A(_8076_), .Y(_6192_) );
OAI21X1 OAI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(_5560_), .B(_5562_), .C(_5555_), .Y(_6193_) );
INVX1 INVX1_819 ( .gnd(gnd), .vdd(vdd), .A(_6193_), .Y(_6194_) );
AND2X2 AND2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_6186_), .B(_6189_), .Y(_6195_) );
AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_8073_), .B(_6192_), .C(_6195_), .D(_6194_), .Y(_6196_) );
NAND3X1 NAND3X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_5953_), .B(_6191_), .C(_6196_), .Y(_6197_) );
INVX1 INVX1_820 ( .gnd(gnd), .vdd(vdd), .A(_5953_), .Y(_6198_) );
NOR2X1 NOR2X1_485 ( .gnd(gnd), .vdd(vdd), .A(_6194_), .B(_6195_), .Y(_6199_) );
NAND2X1 NAND2X1_831 ( .gnd(gnd), .vdd(vdd), .A(_8073_), .B(_6192_), .Y(_6200_) );
OAI21X1 OAI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_6190_), .B(_6193_), .C(_6200_), .Y(_6201_) );
OAI21X1 OAI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(_6199_), .B(_6201_), .C(_6198_), .Y(_6202_) );
AND2X2 AND2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_6197_), .B(_6202_), .Y(_6203_) );
INVX1 INVX1_821 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_151_), .Y(_6204_) );
AOI21X1 AOI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_150_), .B(_5586_), .C(_6204_), .Y(_6205_) );
NOR3X1 NOR3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_5588_), .B(module_1_W_151_), .C(_5591_), .Y(_6206_) );
OAI21X1 OAI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(_6205_), .B(_6206_), .C(_6203_), .Y(_6207_) );
NAND2X1 NAND2X1_832 ( .gnd(gnd), .vdd(vdd), .A(_6202_), .B(_6197_), .Y(_6208_) );
OAI21X1 OAI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(_5591_), .B(_5588_), .C(module_1_W_151_), .Y(_6209_) );
NAND3X1 NAND3X1_1369 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_150_), .B(_6204_), .C(_5586_), .Y(_6210_) );
NAND3X1 NAND3X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_6209_), .B(_6210_), .C(_6208_), .Y(_6211_) );
AND2X2 AND2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_6207_), .B(_6211_), .Y(_6212_) );
OAI21X1 OAI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(_5617_), .B(_5597_), .C(_6212_), .Y(_6213_) );
OAI21X1 OAI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(_5265_), .B(_5618_), .C(_5600_), .Y(_6214_) );
INVX1 INVX1_822 ( .gnd(gnd), .vdd(vdd), .A(_6214_), .Y(_6215_) );
NAND2X1 NAND2X1_833 ( .gnd(gnd), .vdd(vdd), .A(_6211_), .B(_6207_), .Y(_6216_) );
AOI21X1 AOI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(_6216_), .B(_6215_), .C(_8088_), .Y(_6217_) );
NAND3X1 NAND3X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_6027_), .B(_6213_), .C(_6217_), .Y(_6218_) );
NOR2X1 NOR2X1_486 ( .gnd(gnd), .vdd(vdd), .A(_6216_), .B(_6215_), .Y(_6219_) );
INVX1 INVX1_823 ( .gnd(gnd), .vdd(vdd), .A(_8088_), .Y(_6220_) );
OAI21X1 OAI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_6212_), .B(_6214_), .C(_6220_), .Y(_6221_) );
OAI21X1 OAI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(_6221_), .B(_6219_), .C(_5966_), .Y(_6222_) );
NAND2X1 NAND2X1_834 ( .gnd(gnd), .vdd(vdd), .A(_6218_), .B(_6222_), .Y(_6223_) );
AOI21X1 AOI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(_6024_), .B(_6026_), .C(_6223_), .Y(_6224_) );
NAND3X1 NAND3X1_1372 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_166_), .B(module_1_W_167_), .C(_5621_), .Y(_6225_) );
OAI21X1 OAI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_5626_), .B(_5623_), .C(_6025_), .Y(_6226_) );
AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_6218_), .B(_6222_), .C(_6226_), .D(_6225_), .Y(_6227_) );
NOR2X1 NOR2X1_487 ( .gnd(gnd), .vdd(vdd), .A(_6227_), .B(_6224_), .Y(_6228_) );
OAI21X1 OAI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(_5652_), .B(_5632_), .C(_6228_), .Y(_6229_) );
OAI21X1 OAI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_5653_), .B(_5263_), .C(_5635_), .Y(_6230_) );
INVX1 INVX1_824 ( .gnd(gnd), .vdd(vdd), .A(_6230_), .Y(_6231_) );
NAND2X1 NAND2X1_835 ( .gnd(gnd), .vdd(vdd), .A(_6225_), .B(_6226_), .Y(_6232_) );
XNOR2X1 XNOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_6232_), .B(_6223_), .Y(_6233_) );
AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_8096_), .B(_8098_), .C(_6233_), .D(_6231_), .Y(_6234_) );
NAND3X1 NAND3X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_6023_), .B(_6229_), .C(_6234_), .Y(_6235_) );
NOR2X1 NOR2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_6233_), .B(_6231_), .Y(_6236_) );
OAI21X1 OAI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(_6228_), .B(_6230_), .C(_8099_), .Y(_6237_) );
OAI21X1 OAI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_6236_), .B(_6237_), .C(_5976_), .Y(_6238_) );
AND2X2 AND2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_6235_), .B(_6238_), .Y(_6239_) );
INVX1 INVX1_825 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_183_), .Y(_6240_) );
AOI21X1 AOI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_182_), .B(_5656_), .C(_6240_), .Y(_6241_) );
NOR3X1 NOR3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_5658_), .B(module_1_W_183_), .C(_5661_), .Y(_6242_) );
OAI21X1 OAI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(_6241_), .B(_6242_), .C(_6239_), .Y(_6243_) );
NAND2X1 NAND2X1_836 ( .gnd(gnd), .vdd(vdd), .A(_6238_), .B(_6235_), .Y(_6244_) );
OAI21X1 OAI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(_5661_), .B(_5658_), .C(module_1_W_183_), .Y(_6245_) );
NAND3X1 NAND3X1_1374 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_182_), .B(_6240_), .C(_5656_), .Y(_6246_) );
NAND3X1 NAND3X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_6245_), .B(_6246_), .C(_6244_), .Y(_6247_) );
NAND2X1 NAND2X1_837 ( .gnd(gnd), .vdd(vdd), .A(_6247_), .B(_6243_), .Y(_6248_) );
NOR2X1 NOR2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_6248_), .B(_6022_), .Y(_6249_) );
AND2X2 AND2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_6243_), .B(_6247_), .Y(_6250_) );
OAI21X1 OAI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(_6250_), .B(_6021_), .C(_4681_), .Y(_6251_) );
OAI21X1 OAI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(_6251_), .B(_6249_), .C(module_1_W_199_), .Y(_6252_) );
INVX1 INVX1_826 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_199_), .Y(_6253_) );
OAI21X1 OAI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(_5671_), .B(_5690_), .C(_6250_), .Y(_6255_) );
AOI21X1 AOI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(_6248_), .B(_6022_), .C(_8113_), .Y(_6256_) );
NAND3X1 NAND3X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_6253_), .B(_6255_), .C(_6256_), .Y(_6257_) );
NAND2X1 NAND2X1_838 ( .gnd(gnd), .vdd(vdd), .A(_6257_), .B(_6252_), .Y(_6258_) );
NOR3X1 NOR3X1_166 ( .gnd(gnd), .vdd(vdd), .A(_5690_), .B(_5692_), .C(_5691_), .Y(_6259_) );
NOR3X1 NOR3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_5257_), .B(_5697_), .C(_6259_), .Y(_6260_) );
OAI21X1 OAI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(_6260_), .B(_5696_), .C(_5985_), .Y(_6261_) );
INVX2 INVX2_217 ( .gnd(gnd), .vdd(vdd), .A(_5985_), .Y(_6262_) );
NAND3X1 NAND3X1_1377 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_198_), .B(_6262_), .C(_5694_), .Y(_6263_) );
NAND3X1 NAND3X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_6261_), .B(_6263_), .C(_6258_), .Y(_6264_) );
AND2X2 AND2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_6252_), .B(_6257_), .Y(_6266_) );
AOI21X1 AOI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_198_), .B(_5694_), .C(_6262_), .Y(_6267_) );
INVX1 INVX1_827 ( .gnd(gnd), .vdd(vdd), .A(_6263_), .Y(_6268_) );
OAI21X1 OAI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(_6268_), .B(_6267_), .C(_6266_), .Y(_6269_) );
AOI21X1 AOI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(_6264_), .B(_6269_), .C(_6020_), .Y(_6270_) );
OAI21X1 OAI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(_5727_), .B(_5256_), .C(_5707_), .Y(_6271_) );
NAND2X1 NAND2X1_839 ( .gnd(gnd), .vdd(vdd), .A(_6264_), .B(_6269_), .Y(_6272_) );
OAI21X1 OAI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(_6272_), .B(_6271_), .C(_8128_), .Y(_6273_) );
NOR3X1 NOR3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_6270_), .B(_5996_), .C(_6273_), .Y(_6274_) );
INVX2 INVX2_218 ( .gnd(gnd), .vdd(vdd), .A(_5996_), .Y(_6275_) );
INVX1 INVX1_828 ( .gnd(gnd), .vdd(vdd), .A(_6270_), .Y(_6277_) );
AND2X2 AND2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_6269_), .B(_6264_), .Y(_6278_) );
AOI21X1 AOI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(_6020_), .B(_6278_), .C(_8131_), .Y(_6279_) );
AOI21X1 AOI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(_6277_), .B(_6279_), .C(_6275_), .Y(_6280_) );
NOR2X1 NOR2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_6274_), .B(_6280_), .Y(_6281_) );
INVX1 INVX1_829 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_215_), .Y(_6282_) );
AOI21X1 AOI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_214_), .B(_5730_), .C(_6282_), .Y(_6283_) );
NOR3X1 NOR3X1_169 ( .gnd(gnd), .vdd(vdd), .A(_5732_), .B(module_1_W_215_), .C(_5735_), .Y(_6284_) );
OAI21X1 OAI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_6283_), .B(_6284_), .C(_6281_), .Y(_6285_) );
NAND3X1 NAND3X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_6275_), .B(_6277_), .C(_6279_), .Y(_6286_) );
OAI21X1 OAI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_6273_), .B(_6270_), .C(_5996_), .Y(_6288_) );
NAND2X1 NAND2X1_840 ( .gnd(gnd), .vdd(vdd), .A(_6288_), .B(_6286_), .Y(_6289_) );
OAI21X1 OAI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_5735_), .B(_5732_), .C(module_1_W_215_), .Y(_6290_) );
NAND3X1 NAND3X1_1380 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_214_), .B(_6282_), .C(_5730_), .Y(_6291_) );
NAND3X1 NAND3X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_6290_), .B(_6291_), .C(_6289_), .Y(_6292_) );
AND2X2 AND2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_6285_), .B(_6292_), .Y(_6293_) );
OAI21X1 OAI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_5763_), .B(_5741_), .C(_6293_), .Y(_6294_) );
AOI21X1 AOI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_5745_), .B(_5743_), .C(_5763_), .Y(_6295_) );
NAND2X1 NAND2X1_841 ( .gnd(gnd), .vdd(vdd), .A(_6292_), .B(_6285_), .Y(_6296_) );
AOI21X1 AOI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_6295_), .B(_6296_), .C(_8140_), .Y(_6297_) );
NAND3X1 NAND3X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_6019_), .B(_6297_), .C(_6294_), .Y(_6299_) );
NOR2X1 NOR2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_6295_), .B(_6296_), .Y(_6300_) );
INVX1 INVX1_830 ( .gnd(gnd), .vdd(vdd), .A(_8140_), .Y(_6301_) );
OAI21X1 OAI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(_5764_), .B(_5253_), .C(_5744_), .Y(_6302_) );
OAI21X1 OAI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .B(_6302_), .C(_6301_), .Y(_6303_) );
OAI21X1 OAI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_6303_), .B(_6300_), .C(_6006_), .Y(_6304_) );
AND2X2 AND2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_6304_), .B(_6299_), .Y(_6305_) );
INVX1 INVX1_831 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_231_), .Y(_6306_) );
AOI21X1 AOI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_230_), .B(_5767_), .C(_6306_), .Y(_6307_) );
NOR3X1 NOR3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_5769_), .B(module_1_W_231_), .C(_5772_), .Y(_6308_) );
OAI21X1 OAI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(_6307_), .B(_6308_), .C(_6305_), .Y(_6310_) );
NAND2X1 NAND2X1_842 ( .gnd(gnd), .vdd(vdd), .A(_6299_), .B(_6304_), .Y(_6311_) );
OAI21X1 OAI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(_5772_), .B(_5769_), .C(module_1_W_231_), .Y(_6312_) );
NAND3X1 NAND3X1_1383 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_230_), .B(_6306_), .C(_5767_), .Y(_6313_) );
NAND3X1 NAND3X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_6312_), .B(_6313_), .C(_6311_), .Y(_6314_) );
AND2X2 AND2X2_144 ( .gnd(gnd), .vdd(vdd), .A(_6310_), .B(_6314_), .Y(_6315_) );
OAI21X1 OAI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(_5800_), .B(_5778_), .C(_6315_), .Y(_6316_) );
OAI21X1 OAI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(_5801_), .B(_5247_), .C(_5781_), .Y(_6317_) );
INVX1 INVX1_832 ( .gnd(gnd), .vdd(vdd), .A(_6317_), .Y(_6318_) );
NAND2X1 NAND2X1_843 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_6310_), .Y(_6319_) );
AOI21X1 AOI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(_6319_), .B(_6318_), .C(_8153_), .Y(_6321_) );
NAND3X1 NAND3X1_1385 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_247_), .B(_6316_), .C(_6321_), .Y(_6322_) );
INVX2 INVX2_219 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_247_), .Y(_6323_) );
NOR2X1 NOR2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_6319_), .B(_6318_), .Y(_6324_) );
INVX1 INVX1_833 ( .gnd(gnd), .vdd(vdd), .A(_8153_), .Y(_6325_) );
OAI21X1 OAI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(_6315_), .B(_6317_), .C(_6325_), .Y(_6326_) );
OAI21X1 OAI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_6326_), .B(_6324_), .C(_6323_), .Y(_6327_) );
NAND3X1 NAND3X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_6322_), .B(_6327_), .C(_5805_), .Y(_6328_) );
NOR2X1 NOR2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_5806_), .B(_5809_), .Y(_6329_) );
NOR3X1 NOR3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_6324_), .B(_6323_), .C(_6326_), .Y(_6330_) );
AOI21X1 AOI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_6316_), .B(_6321_), .C(module_1_W_247_), .Y(_6332_) );
OAI21X1 OAI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_6330_), .B(_6332_), .C(_6329_), .Y(_6333_) );
NAND3X1 NAND3X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_6018_), .B(_6328_), .C(_6333_), .Y(_6334_) );
NAND3X1 NAND3X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_6323_), .B(_6316_), .C(_6321_), .Y(_6335_) );
OAI21X1 OAI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(_6326_), .B(_6324_), .C(module_1_W_247_), .Y(_6336_) );
AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_246_), .B(_5804_), .C(_6336_), .D(_6335_), .Y(_6337_) );
AOI21X1 AOI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_6322_), .B(_6327_), .C(_5805_), .Y(_6338_) );
OAI21X1 OAI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_6338_), .B(_6337_), .C(_6017_), .Y(_6339_) );
NAND3X1 NAND3X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_6334_), .B(_6339_), .C(_5842_), .Y(_6340_) );
AOI21X1 AOI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_5805_), .B(_5810_), .C(_5222_), .Y(_6341_) );
OAI21X1 OAI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(_6341_), .B(_5245_), .C(_5817_), .Y(_6343_) );
NOR3X1 NOR3X1_172 ( .gnd(gnd), .vdd(vdd), .A(_6337_), .B(_6017_), .C(_6338_), .Y(_6344_) );
AOI21X1 AOI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(_6328_), .B(_6333_), .C(_6018_), .Y(_6345_) );
OAI21X1 OAI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_6344_), .B(_6345_), .C(_6343_), .Y(_6346_) );
NAND2X1 NAND2X1_844 ( .gnd(gnd), .vdd(vdd), .A(_6346_), .B(_6340_), .Y(_6347_) );
NAND2X1 NAND2X1_845 ( .gnd(gnd), .vdd(vdd), .A(_6347_), .B(_5840_), .Y(_6348_) );
OAI21X1 OAI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(_6344_), .B(_6345_), .C(_5842_), .Y(_6349_) );
NAND3X1 NAND3X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_6334_), .B(_6339_), .C(_6343_), .Y(_6350_) );
NAND2X1 NAND2X1_846 ( .gnd(gnd), .vdd(vdd), .A(_6350_), .B(_6349_), .Y(_6351_) );
NAND3X1 NAND3X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_5244_), .B(_6351_), .C(_5837_), .Y(_6352_) );
NAND2X1 NAND2X1_847 ( .gnd(gnd), .vdd(vdd), .A(_6352_), .B(_6348_), .Y(module_1_H_7_) );
NOR2X1 NOR2X1_494 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_248_), .B(_4769_), .Y(_6354_) );
INVX1 INVX1_834 ( .gnd(gnd), .vdd(vdd), .A(_6354_), .Y(_6355_) );
OAI21X1 OAI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_4764_), .B(_4763_), .C(module_1_W_248_), .Y(_6356_) );
NAND2X1 NAND2X1_848 ( .gnd(gnd), .vdd(vdd), .A(_6356_), .B(_6355_), .Y(module_1_H_16_) );
XNOR2X1 XNOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .B(module_1_W_249_), .Y(_6357_) );
INVX1 INVX1_835 ( .gnd(gnd), .vdd(vdd), .A(_6357_), .Y(_6358_) );
OAI21X1 OAI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_248_), .B(_4769_), .C(_6358_), .Y(_6359_) );
INVX2 INVX2_220 ( .gnd(gnd), .vdd(vdd), .A(_6359_), .Y(_6360_) );
NOR2X1 NOR2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_6355_), .B(_6358_), .Y(_6361_) );
NOR2X1 NOR2X1_496 ( .gnd(gnd), .vdd(vdd), .A(_6361_), .B(_6360_), .Y(module_1_H_17_) );
NOR2X1 NOR2X1_497 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_249_), .B(_5239_), .Y(_6363_) );
INVX1 INVX1_836 ( .gnd(gnd), .vdd(vdd), .A(_6363_), .Y(_6364_) );
NAND2X1 NAND2X1_849 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_250_), .B(_5831_), .Y(_6365_) );
OR2X2 OR2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_5831_), .B(module_1_W_250_), .Y(_6366_) );
AOI21X1 AOI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(_6365_), .B(_6366_), .C(_6364_), .Y(_6367_) );
INVX1 INVX1_837 ( .gnd(gnd), .vdd(vdd), .A(_6367_), .Y(_6368_) );
NAND3X1 NAND3X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_6364_), .B(_6365_), .C(_6366_), .Y(_6369_) );
NAND2X1 NAND2X1_850 ( .gnd(gnd), .vdd(vdd), .A(_6369_), .B(_6368_), .Y(_6370_) );
XNOR2X1 XNOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_6370_), .B(_6360_), .Y(module_1_H_18_) );
OAI21X1 OAI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_6367_), .B(_6359_), .C(_6369_), .Y(_6372_) );
NOR2X1 NOR2X1_498 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_250_), .B(_5832_), .Y(_6373_) );
INVX1 INVX1_838 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_251_), .Y(_6374_) );
OAI21X1 OAI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(_6016_), .B(_6013_), .C(_6374_), .Y(_6375_) );
NAND2X1 NAND2X1_851 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_251_), .B(_6017_), .Y(_6376_) );
NAND3X1 NAND3X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_6373_), .B(_6375_), .C(_6376_), .Y(_6377_) );
AOI21X1 AOI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_6375_), .B(_6376_), .C(_6373_), .Y(_6378_) );
INVX1 INVX1_839 ( .gnd(gnd), .vdd(vdd), .A(_6378_), .Y(_6379_) );
NAND2X1 NAND2X1_852 ( .gnd(gnd), .vdd(vdd), .A(_6377_), .B(_6379_), .Y(_6380_) );
XNOR2X1 XNOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_6380_), .B(_6372_), .Y(module_1_H_19_) );
AOI21X1 AOI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_6372_), .B(_6377_), .C(_6378_), .Y(_6382_) );
OAI21X1 OAI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(_5843_), .B(_6011_), .C(_6009_), .Y(_6383_) );
INVX2 INVX2_221 ( .gnd(gnd), .vdd(vdd), .A(_6008_), .Y(_6384_) );
OAI21X1 OAI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_5998_), .B(_5997_), .C(_5788_), .Y(_6385_) );
AOI21X1 AOI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_6385_), .B(_5844_), .C(_5999_), .Y(_6386_) );
NOR3X1 NOR3X1_173 ( .gnd(gnd), .vdd(vdd), .A(_5751_), .B(_5987_), .C(_5990_), .Y(_6387_) );
AOI21X1 AOI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_5991_), .B(_5994_), .C(_6387_), .Y(_6388_) );
OAI21X1 OAI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_5983_), .B(_5980_), .C(_5978_), .Y(_6389_) );
INVX1 INVX1_840 ( .gnd(gnd), .vdd(vdd), .A(_5977_), .Y(_6390_) );
OR2X2 OR2X2_144 ( .gnd(gnd), .vdd(vdd), .A(_5968_), .B(_5851_), .Y(_6391_) );
OAI21X1 OAI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_5970_), .B(_5849_), .C(_6391_), .Y(_6393_) );
NOR2X1 NOR2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_5852_), .B(_6027_), .Y(_6394_) );
OAI21X1 OAI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_5955_), .B(_5956_), .C(_5641_), .Y(_6395_) );
AOI21X1 AOI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_6395_), .B(_5853_), .C(_5957_), .Y(_6396_) );
OAI21X1 OAI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_5951_), .B(_5855_), .C(_5947_), .Y(_6397_) );
INVX2 INVX2_222 ( .gnd(gnd), .vdd(vdd), .A(_6397_), .Y(_6398_) );
NAND2X1 NAND2X1_853 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_139_), .B(_5944_), .Y(_6399_) );
AND2X2 AND2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_5941_), .B(_5937_), .Y(_6400_) );
INVX1 INVX1_841 ( .gnd(gnd), .vdd(vdd), .A(_5938_), .Y(_6401_) );
INVX1 INVX1_842 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf3_), .Y(_6402_) );
XNOR2X1 XNOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_4573_), .B(_6897_), .Y(_6404_) );
NAND2X1 NAND2X1_854 ( .gnd(gnd), .vdd(vdd), .A(_5926_), .B(_5931_), .Y(_6405_) );
XOR2X1 XOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .B(_6425_), .Y(_6406_) );
INVX1 INVX1_843 ( .gnd(gnd), .vdd(vdd), .A(_5860_), .Y(_6407_) );
AOI21X1 AOI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_5914_), .B(_5912_), .C(_5488_), .Y(_6408_) );
OAI21X1 OAI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_6407_), .B(_6408_), .C(_5915_), .Y(_6409_) );
XNOR2X1 XNOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_4522_), .B(_6392_), .Y(_6410_) );
OAI21X1 OAI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_5451_), .B(_4818_), .C(_5454_), .Y(_6411_) );
AOI21X1 AOI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_5905_), .B(_6411_), .C(_5904_), .Y(_6412_) );
INVX1 INVX1_844 ( .gnd(gnd), .vdd(vdd), .A(_5901_), .Y(_6413_) );
INVX1 INVX1_845 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf3_), .Y(_6415_) );
AOI21X1 AOI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(_5898_), .B(_5896_), .C(_5893_), .Y(_6416_) );
NOR2X1 NOR2X1_500 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf0_), .B(_5890_), .Y(_6417_) );
INVX1 INVX1_846 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf2_), .Y(_6418_) );
XNOR2X1 XNOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_8283_), .B(_6331_), .Y(_6419_) );
INVX1 INVX1_847 ( .gnd(gnd), .vdd(vdd), .A(_6419_), .Y(_6420_) );
OAI21X1 OAI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_5884_), .B(_5866_), .C(_5882_), .Y(_6421_) );
XNOR2X1 XNOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_8259_), .B(_6309_), .Y(_6422_) );
INVX1 INVX1_848 ( .gnd(gnd), .vdd(vdd), .A(_6422_), .Y(_6423_) );
AOI21X1 AOI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_5338_), .B(_4796_), .C(_5342_), .Y(_6424_) );
OAI21X1 OAI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_6424_), .B(_5876_), .C(_5874_), .Y(_6426_) );
INVX1 INVX1_849 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_28_), .Y(_6427_) );
XNOR2X1 XNOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_0_), .B(module_1_W_12_), .Y(_6428_) );
XOR2X1 XOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_6428_), .B(module_1_W_8_), .Y(_6429_) );
NAND2X1 NAND2X1_855 ( .gnd(gnd), .vdd(vdd), .A(_6427_), .B(_6429_), .Y(_6430_) );
XNOR2X1 XNOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_6428_), .B(module_1_W_8_), .Y(_6431_) );
NAND2X1 NAND2X1_856 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_28_), .B(_6431_), .Y(_6432_) );
NAND3X1 NAND3X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_5870_), .B(_6432_), .C(_6430_), .Y(_6433_) );
AOI21X1 AOI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_6432_), .B(_6430_), .C(_5870_), .Y(_6434_) );
INVX2 INVX2_223 ( .gnd(gnd), .vdd(vdd), .A(_6434_), .Y(_6435_) );
AOI21X1 AOI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_6433_), .B(_6435_), .C(_6426_), .Y(_6437_) );
INVX1 INVX1_850 ( .gnd(gnd), .vdd(vdd), .A(_5874_), .Y(_6438_) );
AOI21X1 AOI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(_5875_), .B(_5869_), .C(_6438_), .Y(_6439_) );
INVX2 INVX2_224 ( .gnd(gnd), .vdd(vdd), .A(_6433_), .Y(_6440_) );
NOR3X1 NOR3X1_174 ( .gnd(gnd), .vdd(vdd), .A(_6439_), .B(_6434_), .C(_6440_), .Y(_6441_) );
OAI21X1 OAI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_6441_), .B(_6437_), .C(_6423_), .Y(_6442_) );
OAI21X1 OAI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_6440_), .B(_6434_), .C(_6439_), .Y(_6443_) );
NAND3X1 NAND3X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .B(_6433_), .C(_6435_), .Y(_6444_) );
NAND3X1 NAND3X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_6422_), .B(_6444_), .C(_6443_), .Y(_6445_) );
NAND3X1 NAND3X1_1397 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf2_), .B(_6445_), .C(_6442_), .Y(_6446_) );
INVX1 INVX1_851 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf1_), .Y(_6448_) );
NAND3X1 NAND3X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_6423_), .B(_6444_), .C(_6443_), .Y(_6449_) );
OAI21X1 OAI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_6441_), .B(_6437_), .C(_6422_), .Y(_6450_) );
NAND3X1 NAND3X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_6448_), .B(_6449_), .C(_6450_), .Y(_6451_) );
NAND3X1 NAND3X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_5878_), .B(_6446_), .C(_6451_), .Y(_6452_) );
INVX1 INVX1_852 ( .gnd(gnd), .vdd(vdd), .A(_5878_), .Y(_6453_) );
NAND3X1 NAND3X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_6448_), .B(_6445_), .C(_6442_), .Y(_6454_) );
NAND3X1 NAND3X1_1402 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf0_), .B(_6449_), .C(_6450_), .Y(_6455_) );
NAND3X1 NAND3X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_6453_), .B(_6454_), .C(_6455_), .Y(_6456_) );
AOI21X1 AOI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_6452_), .B(_6456_), .C(_6421_), .Y(_6457_) );
INVX1 INVX1_853 ( .gnd(gnd), .vdd(vdd), .A(_5882_), .Y(_6459_) );
AOI21X1 AOI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(_5883_), .B(_5889_), .C(_6459_), .Y(_6460_) );
AOI21X1 AOI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(_6454_), .B(_6455_), .C(_6453_), .Y(_6461_) );
AOI21X1 AOI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_6446_), .B(_6451_), .C(_5878_), .Y(_6462_) );
NOR3X1 NOR3X1_175 ( .gnd(gnd), .vdd(vdd), .A(_6461_), .B(_6460_), .C(_6462_), .Y(_6463_) );
OAI21X1 OAI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_6463_), .B(_6457_), .C(_6420_), .Y(_6464_) );
OAI21X1 OAI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_6461_), .B(_6462_), .C(_6460_), .Y(_6465_) );
NAND3X1 NAND3X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_6452_), .B(_6456_), .C(_6421_), .Y(_6466_) );
NAND3X1 NAND3X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_6419_), .B(_6465_), .C(_6466_), .Y(_6467_) );
NAND3X1 NAND3X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_6418_), .B(_6467_), .C(_6464_), .Y(_6468_) );
NAND3X1 NAND3X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_6420_), .B(_6465_), .C(_6466_), .Y(_6470_) );
OAI21X1 OAI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_6463_), .B(_6457_), .C(_6419_), .Y(_6471_) );
NAND3X1 NAND3X1_1408 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf1_), .B(_6470_), .C(_6471_), .Y(_6472_) );
AOI21X1 AOI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(_6468_), .B(_6472_), .C(_6417_), .Y(_6473_) );
INVX1 INVX1_854 ( .gnd(gnd), .vdd(vdd), .A(_6417_), .Y(_6474_) );
NAND3X1 NAND3X1_1409 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf0_), .B(_6467_), .C(_6464_), .Y(_6475_) );
NAND3X1 NAND3X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_6418_), .B(_6470_), .C(_6471_), .Y(_6476_) );
AOI21X1 AOI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(_6475_), .B(_6476_), .C(_6474_), .Y(_6477_) );
OAI21X1 OAI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_6473_), .B(_6477_), .C(_6416_), .Y(_6478_) );
OAI21X1 OAI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_5864_), .B(_5894_), .C(_5897_), .Y(_6479_) );
NAND3X1 NAND3X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_6474_), .B(_6475_), .C(_6476_), .Y(_6481_) );
NAND3X1 NAND3X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_6417_), .B(_6468_), .C(_6472_), .Y(_6482_) );
NAND3X1 NAND3X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_6481_), .B(_6482_), .C(_6479_), .Y(_6483_) );
XNOR2X1 XNOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_4497_), .B(_6362_), .Y(_6484_) );
NAND3X1 NAND3X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_6484_), .B(_6483_), .C(_6478_), .Y(_6485_) );
AOI21X1 AOI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_6481_), .B(_6482_), .C(_6479_), .Y(_6486_) );
NOR3X1 NOR3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_6473_), .B(_6477_), .C(_6416_), .Y(_6487_) );
INVX1 INVX1_855 ( .gnd(gnd), .vdd(vdd), .A(_6484_), .Y(_6488_) );
OAI21X1 OAI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_6487_), .B(_6486_), .C(_6488_), .Y(_6489_) );
NAND3X1 NAND3X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_6415_), .B(_6485_), .C(_6489_), .Y(_6490_) );
NAND3X1 NAND3X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_6488_), .B(_6483_), .C(_6478_), .Y(_6492_) );
OAI21X1 OAI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_6487_), .B(_6486_), .C(_6484_), .Y(_6493_) );
NAND3X1 NAND3X1_1417 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf2_), .B(_6492_), .C(_6493_), .Y(_6494_) );
AOI21X1 AOI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_6490_), .B(_6494_), .C(_6413_), .Y(_6495_) );
NAND3X1 NAND3X1_1418 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf1_), .B(_6485_), .C(_6489_), .Y(_6496_) );
NAND3X1 NAND3X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_6415_), .B(_6492_), .C(_6493_), .Y(_6497_) );
AOI21X1 AOI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_6496_), .B(_6497_), .C(_5901_), .Y(_6498_) );
OAI21X1 OAI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_6495_), .B(_6498_), .C(_6412_), .Y(_6499_) );
INVX1 INVX1_856 ( .gnd(gnd), .vdd(vdd), .A(_5904_), .Y(_6500_) );
OAI21X1 OAI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_5861_), .B(_5906_), .C(_6500_), .Y(_6501_) );
NAND3X1 NAND3X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_5901_), .B(_6496_), .C(_6497_), .Y(_6503_) );
NAND3X1 NAND3X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_6413_), .B(_6490_), .C(_6494_), .Y(_6504_) );
NAND3X1 NAND3X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_6503_), .B(_6504_), .C(_6501_), .Y(_6505_) );
NAND3X1 NAND3X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_6410_), .B(_6499_), .C(_6505_), .Y(_6506_) );
INVX1 INVX1_857 ( .gnd(gnd), .vdd(vdd), .A(_6410_), .Y(_6507_) );
AOI21X1 AOI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_6503_), .B(_6504_), .C(_6501_), .Y(_6508_) );
NOR3X1 NOR3X1_177 ( .gnd(gnd), .vdd(vdd), .A(_6495_), .B(_6498_), .C(_6412_), .Y(_6509_) );
OAI21X1 OAI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_6509_), .B(_6508_), .C(_6507_), .Y(_6510_) );
NAND3X1 NAND3X1_1424 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf2_), .B(_6506_), .C(_6510_), .Y(_6511_) );
INVX1 INVX1_858 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf1_), .Y(_6512_) );
NAND3X1 NAND3X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_6507_), .B(_6499_), .C(_6505_), .Y(_6514_) );
OAI21X1 OAI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_6509_), .B(_6508_), .C(_6410_), .Y(_6515_) );
NAND3X1 NAND3X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_6512_), .B(_6514_), .C(_6515_), .Y(_6516_) );
NAND3X1 NAND3X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_5916_), .B(_6511_), .C(_6516_), .Y(_6517_) );
INVX1 INVX1_859 ( .gnd(gnd), .vdd(vdd), .A(_5916_), .Y(_6518_) );
NAND3X1 NAND3X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_6512_), .B(_6506_), .C(_6510_), .Y(_6519_) );
NAND3X1 NAND3X1_1429 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf0_), .B(_6514_), .C(_6515_), .Y(_6520_) );
NAND3X1 NAND3X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_6518_), .B(_6519_), .C(_6520_), .Y(_6521_) );
AOI21X1 AOI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_6517_), .B(_6521_), .C(_6409_), .Y(_6522_) );
AOI21X1 AOI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_5917_), .B(_5916_), .C(_5491_), .Y(_6523_) );
AOI21X1 AOI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_5860_), .B(_5918_), .C(_6523_), .Y(_6525_) );
AOI21X1 AOI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_6519_), .B(_6520_), .C(_6518_), .Y(_6526_) );
AOI21X1 AOI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(_6511_), .B(_6516_), .C(_5916_), .Y(_6527_) );
NOR3X1 NOR3X1_178 ( .gnd(gnd), .vdd(vdd), .A(_6526_), .B(_6527_), .C(_6525_), .Y(_6528_) );
OAI21X1 OAI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_6528_), .B(_6522_), .C(_6406_), .Y(_6529_) );
INVX1 INVX1_860 ( .gnd(gnd), .vdd(vdd), .A(_6406_), .Y(_6530_) );
OAI21X1 OAI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_6526_), .B(_6527_), .C(_6525_), .Y(_6531_) );
NAND3X1 NAND3X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_6517_), .B(_6521_), .C(_6409_), .Y(_6532_) );
NAND3X1 NAND3X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_6530_), .B(_6531_), .C(_6532_), .Y(_6533_) );
NAND3X1 NAND3X1_1433 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf3_), .B(_6533_), .C(_6529_), .Y(_6534_) );
INVX1 INVX1_861 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf2_), .Y(_6536_) );
NAND3X1 NAND3X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_6406_), .B(_6531_), .C(_6532_), .Y(_6537_) );
OAI21X1 OAI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_6528_), .B(_6522_), .C(_6530_), .Y(_6538_) );
NAND3X1 NAND3X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_6536_), .B(_6537_), .C(_6538_), .Y(_6539_) );
NAND3X1 NAND3X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_5927_), .B(_6534_), .C(_6539_), .Y(_6540_) );
INVX1 INVX1_862 ( .gnd(gnd), .vdd(vdd), .A(_5927_), .Y(_6541_) );
NAND3X1 NAND3X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_6536_), .B(_6533_), .C(_6529_), .Y(_6542_) );
NAND3X1 NAND3X1_1438 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf1_), .B(_6537_), .C(_6538_), .Y(_6543_) );
NAND3X1 NAND3X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_6541_), .B(_6542_), .C(_6543_), .Y(_6544_) );
AOI21X1 AOI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_6540_), .B(_6544_), .C(_6405_), .Y(_6545_) );
INVX1 INVX1_863 ( .gnd(gnd), .vdd(vdd), .A(_5926_), .Y(_6547_) );
AOI21X1 AOI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(_5929_), .B(_5858_), .C(_6547_), .Y(_6548_) );
AOI21X1 AOI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(_6542_), .B(_6543_), .C(_6541_), .Y(_6549_) );
AOI21X1 AOI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_6534_), .B(_6539_), .C(_5927_), .Y(_6550_) );
NOR3X1 NOR3X1_179 ( .gnd(gnd), .vdd(vdd), .A(_6549_), .B(_6548_), .C(_6550_), .Y(_6551_) );
OAI21X1 OAI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_6551_), .B(_6545_), .C(_6404_), .Y(_6552_) );
INVX1 INVX1_864 ( .gnd(gnd), .vdd(vdd), .A(_6404_), .Y(_6553_) );
OAI21X1 OAI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_6549_), .B(_6550_), .C(_6548_), .Y(_6554_) );
NAND3X1 NAND3X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_6540_), .B(_6544_), .C(_6405_), .Y(_6555_) );
NAND3X1 NAND3X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_6553_), .B(_6555_), .C(_6554_), .Y(_6556_) );
NAND3X1 NAND3X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_6402_), .B(_6556_), .C(_6552_), .Y(_6558_) );
NAND3X1 NAND3X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_6404_), .B(_6555_), .C(_6554_), .Y(_6559_) );
OAI21X1 OAI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_6551_), .B(_6545_), .C(_6553_), .Y(_6560_) );
NAND3X1 NAND3X1_1444 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf2_), .B(_6559_), .C(_6560_), .Y(_6561_) );
AOI21X1 AOI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(_6558_), .B(_6561_), .C(_6401_), .Y(_6562_) );
NAND3X1 NAND3X1_1445 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf1_), .B(_6556_), .C(_6552_), .Y(_6563_) );
NAND3X1 NAND3X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_6402_), .B(_6559_), .C(_6560_), .Y(_6564_) );
AOI21X1 AOI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_6563_), .B(_6564_), .C(_5938_), .Y(_6565_) );
OAI21X1 OAI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_6562_), .B(_6565_), .C(_6400_), .Y(_6566_) );
NAND2X1 NAND2X1_857 ( .gnd(gnd), .vdd(vdd), .A(_5937_), .B(_5941_), .Y(_6567_) );
NAND3X1 NAND3X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_5938_), .B(_6563_), .C(_6564_), .Y(_6569_) );
NAND3X1 NAND3X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_6401_), .B(_6558_), .C(_6561_), .Y(_6570_) );
NAND3X1 NAND3X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_6567_), .B(_6569_), .C(_6570_), .Y(_6571_) );
NAND3X1 NAND3X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_6875_), .B(_6571_), .C(_6566_), .Y(_6572_) );
AOI21X1 AOI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(_6569_), .B(_6570_), .C(_6567_), .Y(_6573_) );
NOR3X1 NOR3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_6565_), .B(_6400_), .C(_6562_), .Y(_6574_) );
OAI21X1 OAI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_6574_), .B(_6573_), .C(_6491_), .Y(_6575_) );
NAND2X1 NAND2X1_858 ( .gnd(gnd), .vdd(vdd), .A(_6572_), .B(_6575_), .Y(_6576_) );
NAND3X1 NAND3X1_1451 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_140_), .B(_4597_), .C(_6576_), .Y(_6577_) );
INVX1 INVX1_865 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_140_), .Y(_6578_) );
OAI21X1 OAI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_6574_), .B(_6573_), .C(_6875_), .Y(_6580_) );
NAND3X1 NAND3X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_6491_), .B(_6571_), .C(_6566_), .Y(_6581_) );
NAND3X1 NAND3X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_4597_), .B(_6581_), .C(_6580_), .Y(_6582_) );
NAND2X1 NAND2X1_859 ( .gnd(gnd), .vdd(vdd), .A(_6578_), .B(_6582_), .Y(_6583_) );
AOI21X1 AOI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(_6577_), .B(_6583_), .C(_6399_), .Y(_6584_) );
INVX1 INVX1_866 ( .gnd(gnd), .vdd(vdd), .A(_6399_), .Y(_6585_) );
NAND2X1 NAND2X1_860 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_140_), .B(_6582_), .Y(_6586_) );
NAND3X1 NAND3X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_6578_), .B(_4597_), .C(_6576_), .Y(_6587_) );
AOI21X1 AOI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_6586_), .B(_6587_), .C(_6585_), .Y(_6588_) );
OAI21X1 OAI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_6588_), .B(_6584_), .C(_6398_), .Y(_6589_) );
NAND3X1 NAND3X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_6585_), .B(_6586_), .C(_6587_), .Y(_6591_) );
NAND3X1 NAND3X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_6399_), .B(_6577_), .C(_6583_), .Y(_6592_) );
NAND3X1 NAND3X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_6397_), .B(_6591_), .C(_6592_), .Y(_6593_) );
NAND3X1 NAND3X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_6524_), .B(_6593_), .C(_6589_), .Y(_6594_) );
NAND2X1 NAND2X1_861 ( .gnd(gnd), .vdd(vdd), .A(_6593_), .B(_6589_), .Y(_6595_) );
AOI21X1 AOI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_6842_), .B(_6595_), .C(_4626_), .Y(_6596_) );
NAND3X1 NAND3X1_1459 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_156_), .B(_6594_), .C(_6596_), .Y(_6597_) );
INVX1 INVX1_867 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_156_), .Y(_6598_) );
AOI21X1 AOI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(_6591_), .B(_6592_), .C(_6397_), .Y(_6599_) );
NOR3X1 NOR3X1_181 ( .gnd(gnd), .vdd(vdd), .A(_6584_), .B(_6588_), .C(_6398_), .Y(_6600_) );
OAI21X1 OAI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_6600_), .B(_6599_), .C(_6842_), .Y(_6602_) );
NAND3X1 NAND3X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_4623_), .B(_6594_), .C(_6602_), .Y(_6603_) );
NAND2X1 NAND2X1_862 ( .gnd(gnd), .vdd(vdd), .A(_6598_), .B(_6603_), .Y(_6604_) );
AOI21X1 AOI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(_6597_), .B(_6604_), .C(_5958_), .Y(_6605_) );
NAND2X1 NAND2X1_863 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_156_), .B(_6603_), .Y(_6606_) );
NAND3X1 NAND3X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_6598_), .B(_6594_), .C(_6596_), .Y(_6607_) );
AOI21X1 AOI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_6607_), .B(_6606_), .C(_5956_), .Y(_6608_) );
OAI21X1 OAI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_6608_), .B(_6605_), .C(_6396_), .Y(_6609_) );
NAND3X1 NAND3X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_5640_), .B(_5954_), .C(_5958_), .Y(_6610_) );
OAI21X1 OAI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_5962_), .B(_5959_), .C(_6610_), .Y(_6611_) );
NAND3X1 NAND3X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_5956_), .B(_6607_), .C(_6606_), .Y(_6613_) );
NAND3X1 NAND3X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_5958_), .B(_6597_), .C(_6604_), .Y(_6614_) );
NAND3X1 NAND3X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_6611_), .B(_6613_), .C(_6614_), .Y(_6615_) );
AOI21X1 AOI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(_6615_), .B(_6609_), .C(_6557_), .Y(_6616_) );
NAND2X1 NAND2X1_864 ( .gnd(gnd), .vdd(vdd), .A(_6615_), .B(_6609_), .Y(_6617_) );
OAI21X1 OAI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_6617_), .B(_6809_), .C(_4648_), .Y(_6618_) );
OAI21X1 OAI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_6618_), .B(_6616_), .C(module_1_W_172_), .Y(_6619_) );
INVX1 INVX1_868 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_172_), .Y(_6620_) );
NAND3X1 NAND3X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_6809_), .B(_6615_), .C(_6609_), .Y(_6621_) );
AOI21X1 AOI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_6613_), .B(_6614_), .C(_6611_), .Y(_6622_) );
NOR3X1 NOR3X1_182 ( .gnd(gnd), .vdd(vdd), .A(_6605_), .B(_6396_), .C(_6608_), .Y(_6624_) );
OAI21X1 OAI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_6624_), .B(_6622_), .C(_6557_), .Y(_6625_) );
NAND2X1 NAND2X1_865 ( .gnd(gnd), .vdd(vdd), .A(_6621_), .B(_6625_), .Y(_6626_) );
NAND3X1 NAND3X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_6620_), .B(_4648_), .C(_6626_), .Y(_6627_) );
NAND3X1 NAND3X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_6394_), .B(_6619_), .C(_6627_), .Y(_6628_) );
NAND3X1 NAND3X1_1469 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_172_), .B(_4648_), .C(_6626_), .Y(_6629_) );
OAI21X1 OAI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_6618_), .B(_6616_), .C(_6620_), .Y(_6630_) );
NAND3X1 NAND3X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_5967_), .B(_6630_), .C(_6629_), .Y(_6631_) );
AOI21X1 AOI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(_6628_), .B(_6631_), .C(_6393_), .Y(_6632_) );
INVX1 INVX1_869 ( .gnd(gnd), .vdd(vdd), .A(_5970_), .Y(_6633_) );
AOI21X1 AOI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(_6633_), .B(_5850_), .C(_5969_), .Y(_6635_) );
AOI21X1 AOI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(_6630_), .B(_6629_), .C(_5967_), .Y(_6636_) );
AOI21X1 AOI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(_6619_), .B(_6627_), .C(_6394_), .Y(_6637_) );
NOR3X1 NOR3X1_183 ( .gnd(gnd), .vdd(vdd), .A(_6636_), .B(_6637_), .C(_6635_), .Y(_6638_) );
OAI21X1 OAI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_6638_), .B(_6632_), .C(_6787_), .Y(_6639_) );
OAI21X1 OAI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_6637_), .B(_6636_), .C(_6635_), .Y(_6640_) );
NAND3X1 NAND3X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_6393_), .B(_6628_), .C(_6631_), .Y(_6641_) );
NAND3X1 NAND3X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_6590_), .B(_6641_), .C(_6640_), .Y(_6642_) );
NAND3X1 NAND3X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_4667_), .B(_6642_), .C(_6639_), .Y(_6643_) );
NAND2X1 NAND2X1_866 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_188_), .B(_6643_), .Y(_6644_) );
INVX1 INVX1_870 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_188_), .Y(_6646_) );
NAND3X1 NAND3X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_6787_), .B(_6641_), .C(_6640_), .Y(_6647_) );
OAI21X1 OAI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_6638_), .B(_6632_), .C(_6590_), .Y(_6648_) );
NAND2X1 NAND2X1_867 ( .gnd(gnd), .vdd(vdd), .A(_6647_), .B(_6648_), .Y(_6649_) );
NAND3X1 NAND3X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_6646_), .B(_4667_), .C(_6649_), .Y(_6650_) );
NAND3X1 NAND3X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_6390_), .B(_6644_), .C(_6650_), .Y(_6651_) );
NAND3X1 NAND3X1_1477 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_188_), .B(_4667_), .C(_6649_), .Y(_6652_) );
NAND2X1 NAND2X1_868 ( .gnd(gnd), .vdd(vdd), .A(_6646_), .B(_6643_), .Y(_6653_) );
NAND3X1 NAND3X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_5977_), .B(_6652_), .C(_6653_), .Y(_6654_) );
AOI21X1 AOI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(_6651_), .B(_6654_), .C(_6389_), .Y(_6655_) );
INVX1 INVX1_871 ( .gnd(gnd), .vdd(vdd), .A(_5980_), .Y(_6657_) );
AOI21X1 AOI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(_5847_), .B(_6657_), .C(_5979_), .Y(_6658_) );
AOI21X1 AOI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(_6652_), .B(_6653_), .C(_5977_), .Y(_6659_) );
AOI21X1 AOI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(_6644_), .B(_6650_), .C(_6390_), .Y(_6660_) );
NOR3X1 NOR3X1_184 ( .gnd(gnd), .vdd(vdd), .A(_6659_), .B(_6660_), .C(_6658_), .Y(_6661_) );
OAI21X1 OAI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_6661_), .B(_6655_), .C(_6623_), .Y(_6662_) );
OAI21X1 OAI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_6660_), .B(_6659_), .C(_6658_), .Y(_6663_) );
NAND3X1 NAND3X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_6389_), .B(_6651_), .C(_6654_), .Y(_6664_) );
NAND3X1 NAND3X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_6754_), .B(_6664_), .C(_6663_), .Y(_6665_) );
NAND2X1 NAND2X1_869 ( .gnd(gnd), .vdd(vdd), .A(_6665_), .B(_6662_), .Y(_6666_) );
NAND3X1 NAND3X1_1481 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_204_), .B(_4694_), .C(_6666_), .Y(_6668_) );
INVX1 INVX1_872 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_204_), .Y(_6669_) );
AOI21X1 AOI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(_6664_), .B(_6663_), .C(_6623_), .Y(_6670_) );
NAND2X1 NAND2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_6664_), .B(_6663_), .Y(_6671_) );
OAI21X1 OAI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_6671_), .B(_6754_), .C(_4694_), .Y(_6672_) );
OAI21X1 OAI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_6672_), .B(_6670_), .C(_6669_), .Y(_6673_) );
AOI21X1 AOI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(_6673_), .B(_6668_), .C(_5988_), .Y(_6674_) );
OAI21X1 OAI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_6672_), .B(_6670_), .C(module_1_W_204_), .Y(_6675_) );
NAND3X1 NAND3X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_6669_), .B(_4694_), .C(_6666_), .Y(_6676_) );
AOI21X1 AOI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(_6675_), .B(_6676_), .C(_5987_), .Y(_6677_) );
OAI21X1 OAI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_6677_), .B(_6674_), .C(_6388_), .Y(_6679_) );
AOI21X1 AOI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(_5986_), .B(_5988_), .C(_5750_), .Y(_6680_) );
OAI21X1 OAI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_6680_), .B(_5845_), .C(_5989_), .Y(_6681_) );
NAND3X1 NAND3X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_5987_), .B(_6675_), .C(_6676_), .Y(_6682_) );
NAND3X1 NAND3X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_5988_), .B(_6673_), .C(_6668_), .Y(_6683_) );
NAND3X1 NAND3X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_6682_), .B(_6683_), .C(_6681_), .Y(_6684_) );
NAND3X1 NAND3X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_6733_), .B(_6684_), .C(_6679_), .Y(_6685_) );
AOI21X1 AOI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_6682_), .B(_6683_), .C(_6681_), .Y(_6686_) );
NOR3X1 NOR3X1_185 ( .gnd(gnd), .vdd(vdd), .A(_6674_), .B(_6388_), .C(_6677_), .Y(_6687_) );
OAI21X1 OAI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_6687_), .B(_6686_), .C(_6656_), .Y(_6688_) );
NAND2X1 NAND2X1_871 ( .gnd(gnd), .vdd(vdd), .A(_6685_), .B(_6688_), .Y(_6690_) );
NAND3X1 NAND3X1_1487 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_220_), .B(_4715_), .C(_6690_), .Y(_6691_) );
INVX1 INVX1_873 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_220_), .Y(_6692_) );
AOI21X1 AOI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(_6684_), .B(_6679_), .C(_6656_), .Y(_6693_) );
NAND2X1 NAND2X1_872 ( .gnd(gnd), .vdd(vdd), .A(_6684_), .B(_6679_), .Y(_6694_) );
OAI21X1 OAI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_6694_), .B(_6733_), .C(_4715_), .Y(_6695_) );
OAI21X1 OAI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_6695_), .B(_6693_), .C(_6692_), .Y(_6696_) );
AOI21X1 AOI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_6696_), .B(_6691_), .C(_6001_), .Y(_6697_) );
OAI21X1 OAI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_6695_), .B(_6693_), .C(module_1_W_220_), .Y(_6698_) );
NAND3X1 NAND3X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_6692_), .B(_4715_), .C(_6690_), .Y(_6699_) );
AOI21X1 AOI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(_6698_), .B(_6699_), .C(_5998_), .Y(_6701_) );
OAI21X1 OAI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_6697_), .B(_6701_), .C(_6386_), .Y(_6702_) );
AOI21X1 AOI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(_5784_), .B(_5792_), .C(_5794_), .Y(_6703_) );
NAND3X1 NAND3X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_5787_), .B(_6001_), .C(_6000_), .Y(_6704_) );
OAI21X1 OAI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_6703_), .B(_6002_), .C(_6704_), .Y(_6705_) );
NAND3X1 NAND3X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_5998_), .B(_6698_), .C(_6699_), .Y(_6706_) );
NAND3X1 NAND3X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_6001_), .B(_6696_), .C(_6691_), .Y(_6707_) );
NAND3X1 NAND3X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_6705_), .B(_6706_), .C(_6707_), .Y(_6708_) );
AOI21X1 AOI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(_6708_), .B(_6702_), .C(_6689_), .Y(_6709_) );
NAND2X1 NAND2X1_873 ( .gnd(gnd), .vdd(vdd), .A(_6708_), .B(_6702_), .Y(_6710_) );
OAI21X1 OAI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_6710_), .B(_6700_), .C(_4741_), .Y(_6712_) );
OAI21X1 OAI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_6712_), .B(_6709_), .C(module_1_W_236_), .Y(_6713_) );
INVX1 INVX1_874 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_236_), .Y(_6714_) );
NAND3X1 NAND3X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_6700_), .B(_6708_), .C(_6702_), .Y(_6715_) );
AOI21X1 AOI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(_6706_), .B(_6707_), .C(_6705_), .Y(_6716_) );
NOR3X1 NOR3X1_186 ( .gnd(gnd), .vdd(vdd), .A(_6697_), .B(_6386_), .C(_6701_), .Y(_6717_) );
OAI21X1 OAI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_6717_), .B(_6716_), .C(_6689_), .Y(_6718_) );
NAND2X1 NAND2X1_874 ( .gnd(gnd), .vdd(vdd), .A(_6715_), .B(_6718_), .Y(_6719_) );
NAND3X1 NAND3X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_6714_), .B(_4741_), .C(_6719_), .Y(_6720_) );
NAND3X1 NAND3X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_6384_), .B(_6713_), .C(_6720_), .Y(_6721_) );
NAND3X1 NAND3X1_1496 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_236_), .B(_4741_), .C(_6719_), .Y(_6723_) );
OAI21X1 OAI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_6712_), .B(_6709_), .C(_6714_), .Y(_6724_) );
NAND3X1 NAND3X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_6008_), .B(_6724_), .C(_6723_), .Y(_6725_) );
AOI21X1 AOI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(_6721_), .B(_6725_), .C(_6383_), .Y(_6726_) );
INVX1 INVX1_875 ( .gnd(gnd), .vdd(vdd), .A(_6011_), .Y(_6727_) );
AOI21X1 AOI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(_6014_), .B(_6727_), .C(_6010_), .Y(_6728_) );
NAND3X1 NAND3X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_6384_), .B(_6724_), .C(_6723_), .Y(_6729_) );
NAND3X1 NAND3X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_6008_), .B(_6713_), .C(_6720_), .Y(_6730_) );
AOI21X1 AOI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(_6729_), .B(_6730_), .C(_6728_), .Y(_6731_) );
OAI21X1 OAI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_6731_), .B(_6726_), .C(_7934_), .Y(_6732_) );
AOI21X1 AOI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_6724_), .B(_6723_), .C(_6008_), .Y(_6734_) );
AOI21X1 AOI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(_6713_), .B(_6720_), .C(_6384_), .Y(_6735_) );
OAI21X1 OAI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_6734_), .B(_6735_), .C(_6728_), .Y(_6736_) );
NAND3X1 NAND3X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_6383_), .B(_6721_), .C(_6725_), .Y(_6737_) );
NAND3X1 NAND3X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_7935_), .B(_6737_), .C(_6736_), .Y(_6738_) );
NAND2X1 NAND2X1_875 ( .gnd(gnd), .vdd(vdd), .A(_6738_), .B(_6732_), .Y(_6739_) );
NAND3X1 NAND3X1_1502 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_252_), .B(_4765_), .C(_6739_), .Y(_6740_) );
INVX1 INVX1_876 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_252_), .Y(_6741_) );
AOI21X1 AOI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_6737_), .B(_6736_), .C(_7934_), .Y(_6742_) );
NAND2X1 NAND2X1_876 ( .gnd(gnd), .vdd(vdd), .A(_6737_), .B(_6736_), .Y(_6743_) );
OAI21X1 OAI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_6743_), .B(_7935_), .C(_4765_), .Y(_6745_) );
OAI21X1 OAI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_6745_), .B(_6742_), .C(_6741_), .Y(_6746_) );
AOI21X1 AOI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(_6746_), .B(_6740_), .C(_6375_), .Y(_6747_) );
INVX1 INVX1_877 ( .gnd(gnd), .vdd(vdd), .A(_6747_), .Y(_6748_) );
NAND3X1 NAND3X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_6375_), .B(_6746_), .C(_6740_), .Y(_6749_) );
NAND2X1 NAND2X1_877 ( .gnd(gnd), .vdd(vdd), .A(_6749_), .B(_6748_), .Y(_6750_) );
XOR2X1 XOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_6750_), .B(_6382_), .Y(module_1_H_20_) );
OAI21X1 OAI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_6747_), .B(_6382_), .C(_6749_), .Y(_6751_) );
NAND2X1 NAND2X1_878 ( .gnd(gnd), .vdd(vdd), .A(_4765_), .B(_6739_), .Y(_6752_) );
NOR2X1 NOR2X1_501 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_252_), .B(_6752_), .Y(_6753_) );
AOI21X1 AOI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_6383_), .B(_6725_), .C(_6734_), .Y(_6755_) );
INVX1 INVX1_878 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_237_), .Y(_6756_) );
OAI21X1 OAI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_6701_), .B(_6386_), .C(_6706_), .Y(_6757_) );
INVX1 INVX1_879 ( .gnd(gnd), .vdd(vdd), .A(_6698_), .Y(_6758_) );
AOI21X1 AOI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_6683_), .B(_6681_), .C(_6674_), .Y(_6759_) );
INVX1 INVX1_880 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_205_), .Y(_6760_) );
OAI21X1 OAI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_6658_), .B(_6660_), .C(_6651_), .Y(_6761_) );
INVX1 INVX1_881 ( .gnd(gnd), .vdd(vdd), .A(_6644_), .Y(_6762_) );
AOI21X1 AOI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(_6393_), .B(_6631_), .C(_6636_), .Y(_6763_) );
INVX1 INVX1_882 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_173_), .Y(_6764_) );
INVX1 INVX1_883 ( .gnd(gnd), .vdd(vdd), .A(_7705_), .Y(_6766_) );
AOI21X1 AOI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(_6611_), .B(_6614_), .C(_6605_), .Y(_6767_) );
INVX1 INVX1_884 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_157_), .Y(_6768_) );
INVX1 INVX1_885 ( .gnd(gnd), .vdd(vdd), .A(_7621_), .Y(_6769_) );
AOI21X1 AOI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(_6397_), .B(_6592_), .C(_6584_), .Y(_6770_) );
INVX1 INVX1_886 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_141_), .Y(_6771_) );
OAI21X1 OAI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_6565_), .B(_6400_), .C(_6569_), .Y(_6772_) );
INVX1 INVX1_887 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf3_), .Y(_6773_) );
AOI21X1 AOI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(_6544_), .B(_6405_), .C(_6549_), .Y(_6774_) );
INVX1 INVX1_888 ( .gnd(gnd), .vdd(vdd), .A(_6542_), .Y(_6775_) );
INVX1 INVX1_889 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf3_), .Y(_6777_) );
AOI21X1 AOI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(_6521_), .B(_6409_), .C(_6526_), .Y(_6778_) );
INVX1 INVX1_890 ( .gnd(gnd), .vdd(vdd), .A(_6519_), .Y(_6779_) );
INVX1 INVX1_891 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf3_), .Y(_6780_) );
AOI21X1 AOI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(_6504_), .B(_6501_), .C(_6495_), .Y(_6781_) );
INVX1 INVX1_892 ( .gnd(gnd), .vdd(vdd), .A(_6490_), .Y(_6782_) );
INVX1 INVX1_893 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf3_), .Y(_6783_) );
OAI21X1 OAI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_6416_), .B(_6477_), .C(_6481_), .Y(_6784_) );
INVX1 INVX1_894 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf2_), .Y(_6785_) );
AOI21X1 AOI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_6456_), .B(_6421_), .C(_6461_), .Y(_6786_) );
INVX1 INVX1_895 ( .gnd(gnd), .vdd(vdd), .A(_6454_), .Y(_6788_) );
INVX1 INVX1_896 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf3_), .Y(_6789_) );
OAI21X1 OAI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_6440_), .B(_6439_), .C(_6435_), .Y(_6790_) );
INVX1 INVX1_897 ( .gnd(gnd), .vdd(vdd), .A(_6430_), .Y(_6791_) );
XOR2X1 XOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_12_), .B(module_1_W_13_), .Y(_6792_) );
INVX1 INVX1_898 ( .gnd(gnd), .vdd(vdd), .A(_6792_), .Y(_6793_) );
OAI21X1 OAI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_7073_), .B(_7084_), .C(module_1_W_9_), .Y(_6794_) );
NAND2X1 NAND2X1_879 ( .gnd(gnd), .vdd(vdd), .A(_4791_), .B(_4934_), .Y(_6795_) );
NAND2X1 NAND2X1_880 ( .gnd(gnd), .vdd(vdd), .A(_6794_), .B(_6795_), .Y(_6796_) );
NAND2X1 NAND2X1_881 ( .gnd(gnd), .vdd(vdd), .A(_6793_), .B(_6796_), .Y(_6797_) );
NAND3X1 NAND3X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_6792_), .B(_6794_), .C(_6795_), .Y(_6799_) );
AOI21X1 AOI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(_6799_), .B(_6797_), .C(module_1_W_29_), .Y(_6800_) );
INVX1 INVX1_899 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_29_), .Y(_6801_) );
NAND2X1 NAND2X1_882 ( .gnd(gnd), .vdd(vdd), .A(_6792_), .B(_6796_), .Y(_6802_) );
NAND3X1 NAND3X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_6793_), .B(_6794_), .C(_6795_), .Y(_6803_) );
AOI21X1 AOI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(_6803_), .B(_6802_), .C(_6801_), .Y(_6804_) );
OAI21X1 OAI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_6804_), .B(_6800_), .C(_6791_), .Y(_6805_) );
NAND3X1 NAND3X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_6801_), .B(_6803_), .C(_6802_), .Y(_6806_) );
NAND3X1 NAND3X1_1507 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_29_), .B(_6799_), .C(_6797_), .Y(_6807_) );
NAND3X1 NAND3X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_6430_), .B(_6807_), .C(_6806_), .Y(_6808_) );
NAND3X1 NAND3X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_6805_), .B(_6808_), .C(_6790_), .Y(_6810_) );
AOI21X1 AOI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(_6433_), .B(_6426_), .C(_6434_), .Y(_6811_) );
AOI21X1 AOI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_6807_), .B(_6806_), .C(_6430_), .Y(_6812_) );
NOR3X1 NOR3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_6800_), .B(_6791_), .C(_6804_), .Y(_6813_) );
OAI21X1 OAI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_6813_), .B(_6812_), .C(_6811_), .Y(_6814_) );
XNOR2X1 XNOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(_7160_), .Y(_6815_) );
INVX1 INVX1_900 ( .gnd(gnd), .vdd(vdd), .A(_6815_), .Y(_6816_) );
NAND3X1 NAND3X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_6814_), .B(_6816_), .C(_6810_), .Y(_6817_) );
NOR3X1 NOR3X1_188 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_6812_), .C(_6813_), .Y(_6818_) );
AOI21X1 AOI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(_6805_), .B(_6808_), .C(_6790_), .Y(_6819_) );
OAI21X1 OAI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_6818_), .B(_6819_), .C(_6815_), .Y(_6821_) );
NAND3X1 NAND3X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_6789_), .B(_6817_), .C(_6821_), .Y(_6822_) );
NAND3X1 NAND3X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_6814_), .B(_6815_), .C(_6810_), .Y(_6823_) );
OAI21X1 OAI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_6818_), .B(_6819_), .C(_6816_), .Y(_6824_) );
NAND3X1 NAND3X1_1513 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf2_), .B(_6823_), .C(_6824_), .Y(_6825_) );
NAND3X1 NAND3X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_6788_), .B(_6822_), .C(_6825_), .Y(_6826_) );
AOI21X1 AOI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(_6823_), .B(_6824_), .C(bloque_datos_13_bF_buf1_), .Y(_6827_) );
AOI21X1 AOI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(_6817_), .B(_6821_), .C(_6789_), .Y(_6828_) );
OAI21X1 OAI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_6827_), .B(_6828_), .C(_6454_), .Y(_6829_) );
NAND3X1 NAND3X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_6826_), .B(_6829_), .C(_6786_), .Y(_6830_) );
OAI21X1 OAI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_6462_), .B(_6460_), .C(_6452_), .Y(_6832_) );
NAND3X1 NAND3X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_6454_), .B(_6822_), .C(_6825_), .Y(_6833_) );
OAI21X1 OAI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_6827_), .B(_6828_), .C(_6788_), .Y(_6834_) );
NAND3X1 NAND3X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_6833_), .B(_6834_), .C(_6832_), .Y(_6835_) );
XNOR2X1 XNOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_4997_), .B(_7204_), .Y(_6836_) );
INVX1 INVX1_901 ( .gnd(gnd), .vdd(vdd), .A(_6836_), .Y(_6837_) );
NAND3X1 NAND3X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_6835_), .B(_6837_), .C(_6830_), .Y(_6838_) );
AOI21X1 AOI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(_6833_), .B(_6834_), .C(_6832_), .Y(_6839_) );
AOI21X1 AOI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(_6826_), .B(_6829_), .C(_6786_), .Y(_6840_) );
OAI21X1 OAI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_6840_), .B(_6839_), .C(_6836_), .Y(_6841_) );
NAND3X1 NAND3X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_6785_), .B(_6838_), .C(_6841_), .Y(_6843_) );
NOR3X1 NOR3X1_189 ( .gnd(gnd), .vdd(vdd), .A(_6839_), .B(_6836_), .C(_6840_), .Y(_6844_) );
AOI21X1 AOI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_6835_), .B(_6830_), .C(_6837_), .Y(_6845_) );
OAI21X1 OAI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_6844_), .B(_6845_), .C(bloque_datos_29_bF_buf1_), .Y(_6846_) );
NAND3X1 NAND3X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_6468_), .B(_6843_), .C(_6846_), .Y(_6847_) );
INVX1 INVX1_902 ( .gnd(gnd), .vdd(vdd), .A(_6468_), .Y(_6848_) );
NOR3X1 NOR3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(bloque_datos_29_bF_buf0_), .C(_6844_), .Y(_6849_) );
AOI21X1 AOI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(_6838_), .B(_6841_), .C(_6785_), .Y(_6850_) );
OAI21X1 OAI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_6849_), .B(_6850_), .C(_6848_), .Y(_6851_) );
AOI21X1 AOI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_6847_), .B(_6851_), .C(_6784_), .Y(_6852_) );
AOI21X1 AOI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(_6482_), .B(_6479_), .C(_6473_), .Y(_6854_) );
NAND3X1 NAND3X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_6848_), .B(_6843_), .C(_6846_), .Y(_6855_) );
OAI21X1 OAI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_6849_), .B(_6850_), .C(_6468_), .Y(_6856_) );
AOI21X1 AOI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_6855_), .B(_6856_), .C(_6854_), .Y(_6857_) );
XNOR2X1 XNOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_4814_), .B(_7259_), .Y(_6858_) );
NOR3X1 NOR3X1_191 ( .gnd(gnd), .vdd(vdd), .A(_6857_), .B(_6858_), .C(_6852_), .Y(_6859_) );
NAND3X1 NAND3X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_6855_), .B(_6854_), .C(_6856_), .Y(_6860_) );
NAND3X1 NAND3X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_6784_), .B(_6847_), .C(_6851_), .Y(_6861_) );
INVX1 INVX1_903 ( .gnd(gnd), .vdd(vdd), .A(_6858_), .Y(_6862_) );
AOI21X1 AOI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(_6860_), .B(_6861_), .C(_6862_), .Y(_6863_) );
OAI21X1 OAI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_6859_), .B(_6863_), .C(_6783_), .Y(_6865_) );
NAND3X1 NAND3X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_6862_), .B(_6860_), .C(_6861_), .Y(_6866_) );
OAI21X1 OAI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_6852_), .B(_6857_), .C(_6858_), .Y(_6867_) );
NAND3X1 NAND3X1_1525 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf2_), .B(_6866_), .C(_6867_), .Y(_6868_) );
NAND3X1 NAND3X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_6782_), .B(_6868_), .C(_6865_), .Y(_6869_) );
AOI21X1 AOI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_6866_), .B(_6867_), .C(bloque_datos_45_bF_buf1_), .Y(_6870_) );
NOR3X1 NOR3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_6863_), .B(_6783_), .C(_6859_), .Y(_6871_) );
OAI21X1 OAI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_6871_), .B(_6870_), .C(_6490_), .Y(_6872_) );
NAND3X1 NAND3X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_6869_), .B(_6872_), .C(_6781_), .Y(_6873_) );
OAI21X1 OAI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_6412_), .B(_6498_), .C(_6503_), .Y(_6874_) );
NAND3X1 NAND3X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_6490_), .B(_6868_), .C(_6865_), .Y(_6876_) );
OAI21X1 OAI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_6871_), .B(_6870_), .C(_6782_), .Y(_6877_) );
NAND3X1 NAND3X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .B(_6874_), .C(_6877_), .Y(_6878_) );
XOR2X1 XOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_4822_), .B(_7336_), .Y(_6879_) );
INVX1 INVX1_904 ( .gnd(gnd), .vdd(vdd), .A(_6879_), .Y(_6880_) );
NAND3X1 NAND3X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_6880_), .B(_6878_), .C(_6873_), .Y(_6881_) );
AOI21X1 AOI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .B(_6877_), .C(_6874_), .Y(_6882_) );
AOI21X1 AOI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(_6869_), .B(_6872_), .C(_6781_), .Y(_6883_) );
OAI21X1 OAI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_6883_), .B(_6882_), .C(_6879_), .Y(_6884_) );
NAND3X1 NAND3X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_6780_), .B(_6881_), .C(_6884_), .Y(_6885_) );
NAND3X1 NAND3X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_6879_), .B(_6878_), .C(_6873_), .Y(_6887_) );
OAI21X1 OAI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_6883_), .B(_6882_), .C(_6880_), .Y(_6888_) );
NAND3X1 NAND3X1_1533 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf2_), .B(_6887_), .C(_6888_), .Y(_6889_) );
NAND3X1 NAND3X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_6779_), .B(_6885_), .C(_6889_), .Y(_6890_) );
AOI21X1 AOI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(_6887_), .B(_6888_), .C(bloque_datos_61_bF_buf1_), .Y(_6891_) );
AOI21X1 AOI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(_6881_), .B(_6884_), .C(_6780_), .Y(_6892_) );
OAI21X1 OAI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_6891_), .B(_6892_), .C(_6519_), .Y(_6893_) );
NAND3X1 NAND3X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_6890_), .B(_6893_), .C(_6778_), .Y(_6894_) );
OAI21X1 OAI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_6525_), .B(_6527_), .C(_6517_), .Y(_6895_) );
NAND3X1 NAND3X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_6519_), .B(_6885_), .C(_6889_), .Y(_6896_) );
OAI21X1 OAI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_6891_), .B(_6892_), .C(_6779_), .Y(_6898_) );
NAND3X1 NAND3X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_6896_), .B(_6895_), .C(_6898_), .Y(_6899_) );
XNOR2X1 XNOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_4827_), .B(_7402_), .Y(_6900_) );
INVX1 INVX1_905 ( .gnd(gnd), .vdd(vdd), .A(_6900_), .Y(_6901_) );
NAND3X1 NAND3X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_6901_), .B(_6899_), .C(_6894_), .Y(_6902_) );
AOI21X1 AOI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(_6896_), .B(_6898_), .C(_6895_), .Y(_6903_) );
AOI21X1 AOI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(_6890_), .B(_6893_), .C(_6778_), .Y(_6904_) );
OAI21X1 OAI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_6903_), .B(_6904_), .C(_6900_), .Y(_6905_) );
NAND3X1 NAND3X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_6777_), .B(_6902_), .C(_6905_), .Y(_6906_) );
NAND3X1 NAND3X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_6900_), .B(_6899_), .C(_6894_), .Y(_6907_) );
OAI21X1 OAI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_6903_), .B(_6904_), .C(_6901_), .Y(_6909_) );
NAND3X1 NAND3X1_1541 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf2_), .B(_6907_), .C(_6909_), .Y(_6910_) );
NAND3X1 NAND3X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_6775_), .B(_6906_), .C(_6910_), .Y(_6911_) );
AOI21X1 AOI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(_6907_), .B(_6909_), .C(bloque_datos_77_bF_buf1_), .Y(_6912_) );
AOI21X1 AOI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(_6902_), .B(_6905_), .C(_6777_), .Y(_6913_) );
OAI21X1 OAI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_6912_), .B(_6913_), .C(_6542_), .Y(_6914_) );
NAND3X1 NAND3X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_6911_), .B(_6914_), .C(_6774_), .Y(_6915_) );
OAI21X1 OAI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_6550_), .B(_6548_), .C(_6540_), .Y(_6916_) );
NAND3X1 NAND3X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_6542_), .B(_6906_), .C(_6910_), .Y(_6917_) );
OAI21X1 OAI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_6912_), .B(_6913_), .C(_6775_), .Y(_6918_) );
NAND3X1 NAND3X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_6917_), .B(_6916_), .C(_6918_), .Y(_6920_) );
XNOR2X1 XNOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_4833_), .B(_7446_), .Y(_6921_) );
INVX1 INVX1_906 ( .gnd(gnd), .vdd(vdd), .A(_6921_), .Y(_6922_) );
NAND3X1 NAND3X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_6922_), .B(_6920_), .C(_6915_), .Y(_6923_) );
AOI21X1 AOI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(_6917_), .B(_6918_), .C(_6916_), .Y(_6924_) );
AOI21X1 AOI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_6911_), .B(_6914_), .C(_6774_), .Y(_6925_) );
OAI21X1 OAI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_6924_), .B(_6925_), .C(_6921_), .Y(_6926_) );
NAND3X1 NAND3X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_6773_), .B(_6923_), .C(_6926_), .Y(_6927_) );
NOR3X1 NOR3X1_193 ( .gnd(gnd), .vdd(vdd), .A(_6924_), .B(_6921_), .C(_6925_), .Y(_6928_) );
AOI21X1 AOI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_6920_), .B(_6915_), .C(_6922_), .Y(_6929_) );
OAI21X1 OAI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_6928_), .B(_6929_), .C(bloque_datos_93_bF_buf2_), .Y(_6931_) );
NAND3X1 NAND3X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_6558_), .B(_6927_), .C(_6931_), .Y(_6932_) );
INVX1 INVX1_907 ( .gnd(gnd), .vdd(vdd), .A(_6558_), .Y(_6933_) );
NOR3X1 NOR3X1_194 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf1_), .B(_6929_), .C(_6928_), .Y(_6934_) );
AOI21X1 AOI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_6923_), .B(_6926_), .C(_6773_), .Y(_6935_) );
OAI21X1 OAI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_6934_), .B(_6935_), .C(_6933_), .Y(_6936_) );
AOI21X1 AOI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_6932_), .B(_6936_), .C(_6772_), .Y(_6937_) );
AOI21X1 AOI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(_6567_), .B(_6570_), .C(_6562_), .Y(_6938_) );
NAND3X1 NAND3X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_6933_), .B(_6927_), .C(_6931_), .Y(_6939_) );
OAI21X1 OAI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_6934_), .B(_6935_), .C(_6558_), .Y(_6940_) );
AOI21X1 AOI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(_6939_), .B(_6940_), .C(_6938_), .Y(_6942_) );
OAI21X1 OAI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_6937_), .B(_6942_), .C(_7544_), .Y(_6943_) );
NAND3X1 NAND3X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_6938_), .B(_6939_), .C(_6940_), .Y(_6944_) );
NAND3X1 NAND3X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_6772_), .B(_6932_), .C(_6936_), .Y(_6945_) );
NAND3X1 NAND3X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_7555_), .B(_6944_), .C(_6945_), .Y(_6946_) );
NAND2X1 NAND2X1_883 ( .gnd(gnd), .vdd(vdd), .A(_6946_), .B(_6943_), .Y(_6947_) );
NAND3X1 NAND3X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_6771_), .B(_4840_), .C(_6947_), .Y(_6948_) );
OAI21X1 OAI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_6937_), .B(_6942_), .C(_7555_), .Y(_6949_) );
NAND3X1 NAND3X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_7544_), .B(_6944_), .C(_6945_), .Y(_6950_) );
NAND3X1 NAND3X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_4840_), .B(_6950_), .C(_6949_), .Y(_6951_) );
NAND2X1 NAND2X1_884 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_141_), .B(_6951_), .Y(_6953_) );
AOI21X1 AOI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .B(_6953_), .C(_6586_), .Y(_6954_) );
INVX1 INVX1_908 ( .gnd(gnd), .vdd(vdd), .A(_6586_), .Y(_6955_) );
NAND3X1 NAND3X1_1556 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_141_), .B(_4840_), .C(_6947_), .Y(_6956_) );
NAND2X1 NAND2X1_885 ( .gnd(gnd), .vdd(vdd), .A(_6771_), .B(_6951_), .Y(_6957_) );
AOI21X1 AOI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(_6956_), .B(_6957_), .C(_6955_), .Y(_6958_) );
OAI21X1 OAI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_6954_), .B(_6958_), .C(_6770_), .Y(_6959_) );
OAI21X1 OAI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_6398_), .B(_6588_), .C(_6591_), .Y(_6960_) );
NAND3X1 NAND3X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_6955_), .B(_6956_), .C(_6957_), .Y(_6961_) );
NAND3X1 NAND3X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_6586_), .B(_6948_), .C(_6953_), .Y(_6962_) );
NAND3X1 NAND3X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_6961_), .B(_6962_), .C(_6960_), .Y(_6964_) );
NAND3X1 NAND3X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_6769_), .B(_6964_), .C(_6959_), .Y(_6965_) );
AOI21X1 AOI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(_6961_), .B(_6962_), .C(_6960_), .Y(_6966_) );
NOR3X1 NOR3X1_195 ( .gnd(gnd), .vdd(vdd), .A(_6954_), .B(_6770_), .C(_6958_), .Y(_6967_) );
OAI21X1 OAI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_6967_), .B(_6966_), .C(_7621_), .Y(_6968_) );
NAND2X1 NAND2X1_886 ( .gnd(gnd), .vdd(vdd), .A(_6965_), .B(_6968_), .Y(_6969_) );
NAND3X1 NAND3X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_6768_), .B(_4848_), .C(_6969_), .Y(_6970_) );
OAI21X1 OAI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_6967_), .B(_6966_), .C(_6769_), .Y(_6971_) );
NAND3X1 NAND3X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_7621_), .B(_6964_), .C(_6959_), .Y(_6972_) );
NAND3X1 NAND3X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_4848_), .B(_6972_), .C(_6971_), .Y(_6973_) );
NAND2X1 NAND2X1_887 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_157_), .B(_6973_), .Y(_6975_) );
AOI21X1 AOI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(_6970_), .B(_6975_), .C(_6606_), .Y(_6976_) );
INVX1 INVX1_909 ( .gnd(gnd), .vdd(vdd), .A(_6606_), .Y(_6977_) );
NAND3X1 NAND3X1_1564 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_157_), .B(_4848_), .C(_6969_), .Y(_6978_) );
NAND2X1 NAND2X1_888 ( .gnd(gnd), .vdd(vdd), .A(_6768_), .B(_6973_), .Y(_6979_) );
AOI21X1 AOI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(_6978_), .B(_6979_), .C(_6977_), .Y(_6980_) );
OAI21X1 OAI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_6976_), .B(_6980_), .C(_6767_), .Y(_6981_) );
OAI21X1 OAI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_6608_), .B(_6396_), .C(_6613_), .Y(_6982_) );
NAND3X1 NAND3X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_6977_), .B(_6978_), .C(_6979_), .Y(_6983_) );
NAND3X1 NAND3X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_6606_), .B(_6970_), .C(_6975_), .Y(_6984_) );
NAND3X1 NAND3X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_6983_), .B(_6984_), .C(_6982_), .Y(_6986_) );
NAND3X1 NAND3X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_6766_), .B(_6986_), .C(_6981_), .Y(_6987_) );
AOI21X1 AOI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(_6983_), .B(_6984_), .C(_6982_), .Y(_6988_) );
NOR3X1 NOR3X1_196 ( .gnd(gnd), .vdd(vdd), .A(_6976_), .B(_6767_), .C(_6980_), .Y(_6989_) );
OAI21X1 OAI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_6989_), .B(_6988_), .C(_7705_), .Y(_6990_) );
NAND2X1 NAND2X1_889 ( .gnd(gnd), .vdd(vdd), .A(_6987_), .B(_6990_), .Y(_6991_) );
NAND3X1 NAND3X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_6764_), .B(_4856_), .C(_6991_), .Y(_6992_) );
OAI21X1 OAI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_6989_), .B(_6988_), .C(_6766_), .Y(_6993_) );
NAND3X1 NAND3X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_7705_), .B(_6986_), .C(_6981_), .Y(_6994_) );
NAND3X1 NAND3X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_4856_), .B(_6994_), .C(_6993_), .Y(_6995_) );
NAND2X1 NAND2X1_890 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_173_), .B(_6995_), .Y(_6997_) );
AOI21X1 AOI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_6992_), .B(_6997_), .C(_6619_), .Y(_6998_) );
INVX1 INVX1_910 ( .gnd(gnd), .vdd(vdd), .A(_6619_), .Y(_6999_) );
NAND3X1 NAND3X1_1572 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_173_), .B(_4856_), .C(_6991_), .Y(_7000_) );
NAND2X1 NAND2X1_891 ( .gnd(gnd), .vdd(vdd), .A(_6764_), .B(_6995_), .Y(_7001_) );
AOI21X1 AOI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_7000_), .B(_7001_), .C(_6999_), .Y(_7002_) );
OAI21X1 OAI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_6998_), .B(_7002_), .C(_6763_), .Y(_7003_) );
OAI21X1 OAI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_6635_), .B(_6637_), .C(_6628_), .Y(_7004_) );
NAND3X1 NAND3X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_6999_), .B(_7000_), .C(_7001_), .Y(_7005_) );
NAND3X1 NAND3X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_6619_), .B(_6992_), .C(_6997_), .Y(_7006_) );
NAND3X1 NAND3X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_7005_), .B(_7006_), .C(_7004_), .Y(_7008_) );
NAND3X1 NAND3X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_7714_), .B(_7008_), .C(_7003_), .Y(_7009_) );
AOI21X1 AOI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(_7005_), .B(_7006_), .C(_7004_), .Y(_7010_) );
NOR3X1 NOR3X1_197 ( .gnd(gnd), .vdd(vdd), .A(_6998_), .B(_6763_), .C(_7002_), .Y(_7011_) );
OAI21X1 OAI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_7011_), .B(_7010_), .C(_7713_), .Y(_7012_) );
NAND2X1 NAND2X1_892 ( .gnd(gnd), .vdd(vdd), .A(_7009_), .B(_7012_), .Y(_7013_) );
NAND3X1 NAND3X1_1577 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_189_), .B(_4864_), .C(_7013_), .Y(_7014_) );
INVX1 INVX1_911 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_189_), .Y(_7015_) );
OAI21X1 OAI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_7011_), .B(_7010_), .C(_7714_), .Y(_7016_) );
NAND3X1 NAND3X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_7713_), .B(_7008_), .C(_7003_), .Y(_7017_) );
NAND3X1 NAND3X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_4864_), .B(_7017_), .C(_7016_), .Y(_7019_) );
NAND2X1 NAND2X1_893 ( .gnd(gnd), .vdd(vdd), .A(_7015_), .B(_7019_), .Y(_7020_) );
NAND3X1 NAND3X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_6762_), .B(_7014_), .C(_7020_), .Y(_7021_) );
NAND3X1 NAND3X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_7015_), .B(_4864_), .C(_7013_), .Y(_7022_) );
NAND2X1 NAND2X1_894 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_189_), .B(_7019_), .Y(_7023_) );
NAND3X1 NAND3X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_6644_), .B(_7022_), .C(_7023_), .Y(_7024_) );
AOI21X1 AOI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_7021_), .B(_7024_), .C(_6761_), .Y(_7025_) );
AOI21X1 AOI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(_6389_), .B(_6654_), .C(_6659_), .Y(_7026_) );
AOI21X1 AOI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_7022_), .B(_7023_), .C(_6644_), .Y(_7027_) );
AOI21X1 AOI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(_7014_), .B(_7020_), .C(_6762_), .Y(_7028_) );
NOR3X1 NOR3X1_198 ( .gnd(gnd), .vdd(vdd), .A(_7027_), .B(_7026_), .C(_7028_), .Y(_7030_) );
OAI21X1 OAI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_7030_), .B(_7025_), .C(_7722_), .Y(_7031_) );
INVX1 INVX1_912 ( .gnd(gnd), .vdd(vdd), .A(_7722_), .Y(_7032_) );
OAI21X1 OAI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_7027_), .B(_7028_), .C(_7026_), .Y(_7033_) );
NAND3X1 NAND3X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_7021_), .B(_7024_), .C(_6761_), .Y(_7034_) );
NAND3X1 NAND3X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_7032_), .B(_7033_), .C(_7034_), .Y(_7035_) );
NAND2X1 NAND2X1_895 ( .gnd(gnd), .vdd(vdd), .A(_7035_), .B(_7031_), .Y(_7036_) );
NAND3X1 NAND3X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_6760_), .B(_4872_), .C(_7036_), .Y(_7037_) );
OAI21X1 OAI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_7030_), .B(_7025_), .C(_7032_), .Y(_7038_) );
NAND3X1 NAND3X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_7722_), .B(_7033_), .C(_7034_), .Y(_7039_) );
NAND3X1 NAND3X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_4872_), .B(_7039_), .C(_7038_), .Y(_7041_) );
NAND2X1 NAND2X1_896 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_205_), .B(_7041_), .Y(_7042_) );
AOI21X1 AOI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_7037_), .B(_7042_), .C(_6675_), .Y(_7043_) );
INVX1 INVX1_913 ( .gnd(gnd), .vdd(vdd), .A(_6675_), .Y(_7044_) );
NAND3X1 NAND3X1_1588 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_205_), .B(_4872_), .C(_7036_), .Y(_7045_) );
NAND2X1 NAND2X1_897 ( .gnd(gnd), .vdd(vdd), .A(_6760_), .B(_7041_), .Y(_7046_) );
AOI21X1 AOI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(_7045_), .B(_7046_), .C(_7044_), .Y(_7047_) );
OAI21X1 OAI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_7043_), .B(_7047_), .C(_6759_), .Y(_7048_) );
OAI21X1 OAI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_6677_), .B(_6388_), .C(_6682_), .Y(_7049_) );
NAND3X1 NAND3X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_7044_), .B(_7045_), .C(_7046_), .Y(_7050_) );
NAND3X1 NAND3X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_6675_), .B(_7037_), .C(_7042_), .Y(_7052_) );
NAND3X1 NAND3X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_7050_), .B(_7052_), .C(_7049_), .Y(_7053_) );
NAND3X1 NAND3X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_7730_), .B(_7053_), .C(_7048_), .Y(_7054_) );
NAND2X1 NAND2X1_898 ( .gnd(gnd), .vdd(vdd), .A(_7053_), .B(_7048_), .Y(_7055_) );
AOI21X1 AOI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_7731_), .B(_7055_), .C(_4881_), .Y(_7056_) );
NAND3X1 NAND3X1_1593 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_221_), .B(_7054_), .C(_7056_), .Y(_7057_) );
INVX1 INVX1_914 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_221_), .Y(_7058_) );
AOI21X1 AOI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(_7050_), .B(_7052_), .C(_7049_), .Y(_7059_) );
NOR3X1 NOR3X1_199 ( .gnd(gnd), .vdd(vdd), .A(_6759_), .B(_7043_), .C(_7047_), .Y(_7060_) );
OAI21X1 OAI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_7060_), .B(_7059_), .C(_7731_), .Y(_7061_) );
NAND3X1 NAND3X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_4880_), .B(_7054_), .C(_7061_), .Y(_7063_) );
NAND2X1 NAND2X1_899 ( .gnd(gnd), .vdd(vdd), .A(_7058_), .B(_7063_), .Y(_7064_) );
NAND3X1 NAND3X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_6758_), .B(_7057_), .C(_7064_), .Y(_7065_) );
NAND3X1 NAND3X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_7058_), .B(_7054_), .C(_7056_), .Y(_7066_) );
NAND2X1 NAND2X1_900 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_221_), .B(_7063_), .Y(_7067_) );
NAND3X1 NAND3X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_6698_), .B(_7066_), .C(_7067_), .Y(_7068_) );
AOI21X1 AOI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(_7065_), .B(_7068_), .C(_6757_), .Y(_7069_) );
AOI21X1 AOI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_6705_), .B(_6707_), .C(_6697_), .Y(_7070_) );
AOI21X1 AOI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_7066_), .B(_7067_), .C(_6698_), .Y(_7071_) );
AOI21X1 AOI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_7057_), .B(_7064_), .C(_6758_), .Y(_7072_) );
NOR3X1 NOR3X1_200 ( .gnd(gnd), .vdd(vdd), .A(_7071_), .B(_7070_), .C(_7072_), .Y(_7074_) );
OAI21X1 OAI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_7074_), .B(_7069_), .C(_7739_), .Y(_7075_) );
INVX1 INVX1_915 ( .gnd(gnd), .vdd(vdd), .A(_7739_), .Y(_7076_) );
OAI21X1 OAI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_7071_), .B(_7072_), .C(_7070_), .Y(_7077_) );
NAND3X1 NAND3X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_7065_), .B(_7068_), .C(_6757_), .Y(_7078_) );
NAND3X1 NAND3X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_7076_), .B(_7078_), .C(_7077_), .Y(_7079_) );
NAND2X1 NAND2X1_901 ( .gnd(gnd), .vdd(vdd), .A(_7079_), .B(_7075_), .Y(_7080_) );
NAND3X1 NAND3X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_4888_), .C(_7080_), .Y(_7081_) );
OAI21X1 OAI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_7074_), .B(_7069_), .C(_7076_), .Y(_7082_) );
NAND3X1 NAND3X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_7739_), .B(_7078_), .C(_7077_), .Y(_7083_) );
NAND3X1 NAND3X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_7083_), .C(_7082_), .Y(_7085_) );
NAND2X1 NAND2X1_902 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_237_), .B(_7085_), .Y(_7086_) );
AOI21X1 AOI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_7081_), .B(_7086_), .C(_6713_), .Y(_7087_) );
INVX1 INVX1_916 ( .gnd(gnd), .vdd(vdd), .A(_6713_), .Y(_7088_) );
NAND3X1 NAND3X1_1603 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_237_), .B(_4888_), .C(_7080_), .Y(_7089_) );
NAND2X1 NAND2X1_903 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_7085_), .Y(_7090_) );
AOI21X1 AOI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_7089_), .B(_7090_), .C(_7088_), .Y(_7091_) );
OAI21X1 OAI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_7087_), .B(_7091_), .C(_6755_), .Y(_7092_) );
OAI21X1 OAI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_6728_), .B(_6735_), .C(_6721_), .Y(_7093_) );
NAND3X1 NAND3X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_7088_), .B(_7089_), .C(_7090_), .Y(_7094_) );
NAND3X1 NAND3X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_6713_), .B(_7081_), .C(_7086_), .Y(_7096_) );
NAND3X1 NAND3X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_7094_), .B(_7096_), .C(_7093_), .Y(_7097_) );
NAND3X1 NAND3X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_7936_), .B(_7092_), .C(_7097_), .Y(_7098_) );
AOI21X1 AOI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_7094_), .B(_7096_), .C(_7093_), .Y(_7099_) );
NOR3X1 NOR3X1_201 ( .gnd(gnd), .vdd(vdd), .A(_7087_), .B(_6755_), .C(_7091_), .Y(_7100_) );
OAI21X1 OAI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_7100_), .B(_7099_), .C(_7747_), .Y(_7101_) );
NAND2X1 NAND2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_7098_), .B(_7101_), .Y(_7102_) );
NAND3X1 NAND3X1_1608 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_253_), .B(_4896_), .C(_7102_), .Y(_7103_) );
INVX1 INVX1_917 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_253_), .Y(_7104_) );
OAI21X1 OAI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_7100_), .B(_7099_), .C(_7936_), .Y(_7105_) );
NAND3X1 NAND3X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_7747_), .B(_7092_), .C(_7097_), .Y(_7107_) );
NAND3X1 NAND3X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .B(_7107_), .C(_7105_), .Y(_7108_) );
NAND2X1 NAND2X1_905 ( .gnd(gnd), .vdd(vdd), .A(_7104_), .B(_7108_), .Y(_7109_) );
NAND3X1 NAND3X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_6753_), .B(_7103_), .C(_7109_), .Y(_7110_) );
INVX1 INVX1_918 ( .gnd(gnd), .vdd(vdd), .A(_6753_), .Y(_7111_) );
NAND2X1 NAND2X1_906 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_253_), .B(_7108_), .Y(_7112_) );
OR2X2 OR2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_7108_), .B(module_1_W_253_), .Y(_7113_) );
NAND3X1 NAND3X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_7111_), .B(_7112_), .C(_7113_), .Y(_7114_) );
NAND2X1 NAND2X1_907 ( .gnd(gnd), .vdd(vdd), .A(_7110_), .B(_7114_), .Y(_7115_) );
XNOR2X1 XNOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_7115_), .B(_6751_), .Y(module_1_H_21_) );
AOI21X1 AOI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_7103_), .B(_7109_), .C(_6753_), .Y(_7117_) );
AOI21X1 AOI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_6751_), .B(_7110_), .C(_7117_), .Y(_7118_) );
INVX1 INVX1_919 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7119_) );
INVX1 INVX1_920 ( .gnd(gnd), .vdd(vdd), .A(_7112_), .Y(_7120_) );
OAI21X1 OAI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_7091_), .B(_6755_), .C(_7094_), .Y(_7121_) );
OAI21X1 OAI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_7072_), .B(_7070_), .C(_7065_), .Y(_7122_) );
OAI21X1 OAI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_6759_), .B(_7047_), .C(_7050_), .Y(_7123_) );
OAI21X1 OAI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_7028_), .B(_7026_), .C(_7021_), .Y(_7124_) );
INVX1 INVX1_921 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .Y(_7125_) );
INVX1 INVX1_922 ( .gnd(gnd), .vdd(vdd), .A(_7022_), .Y(_7126_) );
OAI21X1 OAI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_7002_), .B(_6763_), .C(_7005_), .Y(_7128_) );
INVX1 INVX1_923 ( .gnd(gnd), .vdd(vdd), .A(_7128_), .Y(_7129_) );
INVX1 INVX1_924 ( .gnd(gnd), .vdd(vdd), .A(_6992_), .Y(_7130_) );
OAI21X1 OAI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_6980_), .B(_6767_), .C(_6983_), .Y(_7131_) );
INVX1 INVX1_925 ( .gnd(gnd), .vdd(vdd), .A(_7131_), .Y(_7132_) );
INVX1 INVX1_926 ( .gnd(gnd), .vdd(vdd), .A(_6970_), .Y(_7133_) );
OAI21X1 OAI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_6958_), .B(_6770_), .C(_6961_), .Y(_7134_) );
NAND2X1 NAND2X1_908 ( .gnd(gnd), .vdd(vdd), .A(_6932_), .B(_6945_), .Y(_7135_) );
INVX1 INVX1_927 ( .gnd(gnd), .vdd(vdd), .A(_7135_), .Y(_7136_) );
NAND2X1 NAND2X1_909 ( .gnd(gnd), .vdd(vdd), .A(_6917_), .B(_6920_), .Y(_7137_) );
NAND2X1 NAND2X1_910 ( .gnd(gnd), .vdd(vdd), .A(_6896_), .B(_6899_), .Y(_7139_) );
NAND2X1 NAND2X1_911 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .B(_6878_), .Y(_7140_) );
NAND2X1 NAND2X1_912 ( .gnd(gnd), .vdd(vdd), .A(_6847_), .B(_6861_), .Y(_7141_) );
NAND2X1 NAND2X1_913 ( .gnd(gnd), .vdd(vdd), .A(_6833_), .B(_6835_), .Y(_7142_) );
OAI21X1 OAI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_6812_), .C(_6808_), .Y(_7143_) );
INVX1 INVX1_928 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_30_), .Y(_7144_) );
NOR2X1 NOR2X1_502 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_12_), .B(module_1_W_13_), .Y(_7145_) );
XNOR2X1 XNOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_7145_), .B(module_1_W_14_), .Y(_7146_) );
XNOR2X1 XNOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_5286_), .B(module_1_W_10_), .Y(_7147_) );
XNOR2X1 XNOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_7147_), .B(_7146_), .Y(_7148_) );
OR2X2 OR2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_7148_), .B(_7144_), .Y(_7150_) );
NAND2X1 NAND2X1_914 ( .gnd(gnd), .vdd(vdd), .A(_7144_), .B(_7148_), .Y(_7151_) );
NAND2X1 NAND2X1_915 ( .gnd(gnd), .vdd(vdd), .A(_7151_), .B(_7150_), .Y(_7152_) );
XNOR2X1 XNOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_7152_), .B(_6804_), .Y(_7153_) );
XOR2X1 XOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_7153_), .B(_7143_), .Y(_7154_) );
XNOR2X1 XNOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_5310_), .B(_5345_), .Y(_7155_) );
XOR2X1 XOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_7154_), .B(_7155_), .Y(_7156_) );
NAND2X1 NAND2X1_916 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf3_), .B(_7156_), .Y(_7157_) );
INVX1 INVX1_929 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf2_), .Y(_7158_) );
XNOR2X1 XNOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_7154_), .B(_7155_), .Y(_7159_) );
NAND2X1 NAND2X1_917 ( .gnd(gnd), .vdd(vdd), .A(_7158_), .B(_7159_), .Y(_7161_) );
NAND3X1 NAND3X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_6828_), .B(_7161_), .C(_7157_), .Y(_7162_) );
NAND2X1 NAND2X1_918 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf1_), .B(_7159_), .Y(_7163_) );
NAND2X1 NAND2X1_919 ( .gnd(gnd), .vdd(vdd), .A(_7158_), .B(_7156_), .Y(_7164_) );
NAND3X1 NAND3X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_6825_), .B(_7163_), .C(_7164_), .Y(_7165_) );
NAND3X1 NAND3X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_7142_), .B(_7162_), .C(_7165_), .Y(_7166_) );
AOI21X1 AOI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_7162_), .B(_7165_), .C(_7142_), .Y(_7167_) );
INVX1 INVX1_930 ( .gnd(gnd), .vdd(vdd), .A(_7167_), .Y(_7168_) );
XNOR2X1 XNOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_5380_), .B(_5331_), .Y(_7169_) );
NAND3X1 NAND3X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_7166_), .B(_7169_), .C(_7168_), .Y(_7170_) );
INVX1 INVX1_931 ( .gnd(gnd), .vdd(vdd), .A(_7166_), .Y(_7172_) );
INVX1 INVX1_932 ( .gnd(gnd), .vdd(vdd), .A(_7169_), .Y(_7173_) );
OAI21X1 OAI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_7172_), .B(_7167_), .C(_7173_), .Y(_7174_) );
NAND3X1 NAND3X1_1617 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf2_), .B(_7170_), .C(_7174_), .Y(_7175_) );
INVX1 INVX1_933 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf1_), .Y(_7176_) );
OAI21X1 OAI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_7172_), .B(_7167_), .C(_7169_), .Y(_7177_) );
NAND3X1 NAND3X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_7166_), .B(_7173_), .C(_7168_), .Y(_7178_) );
NAND3X1 NAND3X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_7176_), .B(_7178_), .C(_7177_), .Y(_7179_) );
NAND3X1 NAND3X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_6850_), .B(_7175_), .C(_7179_), .Y(_7180_) );
NAND3X1 NAND3X1_1621 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf0_), .B(_7178_), .C(_7177_), .Y(_7181_) );
NAND3X1 NAND3X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_7176_), .B(_7170_), .C(_7174_), .Y(_7183_) );
NAND3X1 NAND3X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_6846_), .B(_7181_), .C(_7183_), .Y(_7184_) );
NAND3X1 NAND3X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_7141_), .B(_7180_), .C(_7184_), .Y(_7185_) );
INVX1 INVX1_934 ( .gnd(gnd), .vdd(vdd), .A(_7141_), .Y(_7186_) );
NAND3X1 NAND3X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_6850_), .B(_7181_), .C(_7183_), .Y(_7187_) );
NAND3X1 NAND3X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_6846_), .B(_7175_), .C(_7179_), .Y(_7188_) );
NAND3X1 NAND3X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_7186_), .B(_7187_), .C(_7188_), .Y(_7189_) );
XNOR2X1 XNOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_5418_), .B(_5368_), .Y(_7190_) );
NAND3X1 NAND3X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_7190_), .B(_7185_), .C(_7189_), .Y(_7191_) );
AOI21X1 AOI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_7187_), .B(_7188_), .C(_7186_), .Y(_7192_) );
AOI21X1 AOI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_7180_), .B(_7184_), .C(_7141_), .Y(_7194_) );
INVX1 INVX1_935 ( .gnd(gnd), .vdd(vdd), .A(_7190_), .Y(_7195_) );
OAI21X1 OAI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_7192_), .B(_7194_), .C(_7195_), .Y(_7196_) );
NAND3X1 NAND3X1_1629 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf3_), .B(_7191_), .C(_7196_), .Y(_7197_) );
INVX1 INVX1_936 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf2_), .Y(_7198_) );
OAI21X1 OAI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_7192_), .B(_7194_), .C(_7190_), .Y(_7199_) );
NAND3X1 NAND3X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_7195_), .B(_7185_), .C(_7189_), .Y(_7200_) );
NAND3X1 NAND3X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_7198_), .B(_7200_), .C(_7199_), .Y(_7201_) );
NAND3X1 NAND3X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_6871_), .B(_7197_), .C(_7201_), .Y(_7202_) );
NAND3X1 NAND3X1_1633 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf1_), .B(_7200_), .C(_7199_), .Y(_7203_) );
NAND3X1 NAND3X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_7198_), .B(_7191_), .C(_7196_), .Y(_7205_) );
NAND3X1 NAND3X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_6868_), .B(_7203_), .C(_7205_), .Y(_7206_) );
NAND3X1 NAND3X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_7140_), .B(_7202_), .C(_7206_), .Y(_7207_) );
INVX1 INVX1_937 ( .gnd(gnd), .vdd(vdd), .A(_7140_), .Y(_7208_) );
NAND3X1 NAND3X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_6871_), .B(_7203_), .C(_7205_), .Y(_7209_) );
NAND3X1 NAND3X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_6868_), .B(_7197_), .C(_7201_), .Y(_7210_) );
NAND3X1 NAND3X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_7208_), .B(_7209_), .C(_7210_), .Y(_7211_) );
XNOR2X1 XNOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_5457_), .B(_8034_), .Y(_7212_) );
NAND3X1 NAND3X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_7212_), .B(_7207_), .C(_7211_), .Y(_7213_) );
AOI21X1 AOI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_7209_), .B(_7210_), .C(_7208_), .Y(_7214_) );
AOI21X1 AOI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_7202_), .B(_7206_), .C(_7140_), .Y(_7216_) );
INVX1 INVX1_938 ( .gnd(gnd), .vdd(vdd), .A(_7212_), .Y(_7217_) );
OAI21X1 OAI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_7214_), .B(_7216_), .C(_7217_), .Y(_7218_) );
NAND3X1 NAND3X1_1641 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf2_), .B(_7213_), .C(_7218_), .Y(_7219_) );
INVX1 INVX1_939 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf1_), .Y(_7220_) );
OAI21X1 OAI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_7214_), .B(_7216_), .C(_7212_), .Y(_7221_) );
NAND3X1 NAND3X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_7217_), .B(_7207_), .C(_7211_), .Y(_7222_) );
NAND3X1 NAND3X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_7220_), .B(_7222_), .C(_7221_), .Y(_7223_) );
NAND3X1 NAND3X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_6892_), .B(_7219_), .C(_7223_), .Y(_7224_) );
NAND3X1 NAND3X1_1645 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf0_), .B(_7222_), .C(_7221_), .Y(_7225_) );
NAND3X1 NAND3X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_7220_), .B(_7213_), .C(_7218_), .Y(_7227_) );
NAND3X1 NAND3X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_6889_), .B(_7225_), .C(_7227_), .Y(_7228_) );
NAND3X1 NAND3X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_7139_), .B(_7224_), .C(_7228_), .Y(_7229_) );
INVX2 INVX2_225 ( .gnd(gnd), .vdd(vdd), .A(_7139_), .Y(_7230_) );
AOI21X1 AOI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_7225_), .B(_7227_), .C(_6889_), .Y(_7231_) );
AOI21X1 AOI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_7219_), .B(_7223_), .C(_6892_), .Y(_7232_) );
OAI21X1 OAI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_7231_), .B(_7232_), .C(_7230_), .Y(_7233_) );
XOR2X1 XOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_5498_), .B(_5459_), .Y(_7234_) );
NAND3X1 NAND3X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_7229_), .B(_7234_), .C(_7233_), .Y(_7235_) );
NOR3X1 NOR3X1_202 ( .gnd(gnd), .vdd(vdd), .A(_7231_), .B(_7230_), .C(_7232_), .Y(_7236_) );
AOI21X1 AOI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_7224_), .B(_7228_), .C(_7139_), .Y(_7238_) );
INVX1 INVX1_940 ( .gnd(gnd), .vdd(vdd), .A(_7234_), .Y(_7239_) );
OAI21X1 OAI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_7236_), .B(_7238_), .C(_7239_), .Y(_7240_) );
NAND3X1 NAND3X1_1650 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf3_), .B(_7235_), .C(_7240_), .Y(_7241_) );
INVX1 INVX1_941 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf2_), .Y(_7242_) );
OAI21X1 OAI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_7236_), .B(_7238_), .C(_7234_), .Y(_7243_) );
NAND3X1 NAND3X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_7229_), .B(_7239_), .C(_7233_), .Y(_7244_) );
NAND3X1 NAND3X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_7242_), .B(_7244_), .C(_7243_), .Y(_7245_) );
NAND3X1 NAND3X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_6913_), .B(_7241_), .C(_7245_), .Y(_7246_) );
NAND3X1 NAND3X1_1654 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf1_), .B(_7244_), .C(_7243_), .Y(_7247_) );
NAND3X1 NAND3X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_7242_), .B(_7235_), .C(_7240_), .Y(_7249_) );
NAND3X1 NAND3X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_6910_), .B(_7247_), .C(_7249_), .Y(_7250_) );
NAND3X1 NAND3X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_7137_), .B(_7246_), .C(_7250_), .Y(_7251_) );
INVX1 INVX1_942 ( .gnd(gnd), .vdd(vdd), .A(_7137_), .Y(_7252_) );
NAND3X1 NAND3X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_6913_), .B(_7247_), .C(_7249_), .Y(_7253_) );
NAND3X1 NAND3X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_6910_), .B(_7241_), .C(_7245_), .Y(_7254_) );
NAND3X1 NAND3X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_7252_), .B(_7253_), .C(_7254_), .Y(_7255_) );
XOR2X1 XOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_5538_), .B(_5500_), .Y(_7256_) );
INVX1 INVX1_943 ( .gnd(gnd), .vdd(vdd), .A(_7256_), .Y(_7257_) );
NAND3X1 NAND3X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_7257_), .B(_7251_), .C(_7255_), .Y(_7258_) );
AOI21X1 AOI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_7253_), .B(_7254_), .C(_7252_), .Y(_7260_) );
AOI21X1 AOI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_7246_), .B(_7250_), .C(_7137_), .Y(_7261_) );
OAI21X1 OAI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(_7261_), .C(_7256_), .Y(_7262_) );
NAND3X1 NAND3X1_1662 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf3_), .B(_7258_), .C(_7262_), .Y(_7263_) );
INVX1 INVX1_944 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf2_), .Y(_7264_) );
NAND3X1 NAND3X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_7256_), .B(_7251_), .C(_7255_), .Y(_7265_) );
OAI21X1 OAI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(_7261_), .C(_7257_), .Y(_7266_) );
NAND3X1 NAND3X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_7264_), .B(_7265_), .C(_7266_), .Y(_7267_) );
NAND3X1 NAND3X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_6935_), .B(_7263_), .C(_7267_), .Y(_7268_) );
NAND3X1 NAND3X1_1666 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf1_), .B(_7265_), .C(_7266_), .Y(_7269_) );
NAND3X1 NAND3X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_7264_), .B(_7258_), .C(_7262_), .Y(_7271_) );
NAND3X1 NAND3X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_6931_), .B(_7269_), .C(_7271_), .Y(_7272_) );
AOI21X1 AOI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_7268_), .B(_7272_), .C(_7136_), .Y(_7273_) );
NAND3X1 NAND3X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_6935_), .B(_7269_), .C(_7271_), .Y(_7274_) );
NAND3X1 NAND3X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_6931_), .B(_7263_), .C(_7267_), .Y(_7275_) );
AOI21X1 AOI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_7274_), .B(_7275_), .C(_7135_), .Y(_7276_) );
OAI21X1 OAI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_7273_), .B(_7276_), .C(_5540_), .Y(_7277_) );
INVX1 INVX1_945 ( .gnd(gnd), .vdd(vdd), .A(_5540_), .Y(_7278_) );
NAND3X1 NAND3X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_7135_), .B(_7274_), .C(_7275_), .Y(_7279_) );
NAND3X1 NAND3X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_7268_), .B(_7272_), .C(_7136_), .Y(_7280_) );
NAND3X1 NAND3X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_7278_), .B(_7279_), .C(_7280_), .Y(_7282_) );
NAND3X1 NAND3X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_5579_), .B(_7282_), .C(_7277_), .Y(_7283_) );
NAND2X1 NAND2X1_920 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_142_), .B(_7283_), .Y(_7284_) );
INVX1 INVX1_946 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_142_), .Y(_7285_) );
OAI21X1 OAI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_7273_), .B(_7276_), .C(_7278_), .Y(_7286_) );
NAND3X1 NAND3X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_5540_), .B(_7279_), .C(_7280_), .Y(_7287_) );
NAND2X1 NAND2X1_921 ( .gnd(gnd), .vdd(vdd), .A(_7287_), .B(_7286_), .Y(_7288_) );
NAND3X1 NAND3X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_7285_), .B(_5579_), .C(_7288_), .Y(_7289_) );
NAND3X1 NAND3X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .B(_7289_), .C(_7284_), .Y(_7290_) );
INVX1 INVX1_947 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .Y(_7291_) );
NAND3X1 NAND3X1_1678 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_142_), .B(_5579_), .C(_7288_), .Y(_7293_) );
NAND2X1 NAND2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_7285_), .B(_7283_), .Y(_7294_) );
NAND3X1 NAND3X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_7291_), .B(_7293_), .C(_7294_), .Y(_7295_) );
NAND3X1 NAND3X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_7134_), .B(_7290_), .C(_7295_), .Y(_7296_) );
INVX1 INVX1_948 ( .gnd(gnd), .vdd(vdd), .A(_7134_), .Y(_7297_) );
NAND3X1 NAND3X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_7291_), .B(_7289_), .C(_7284_), .Y(_7298_) );
NAND3X1 NAND3X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .B(_7293_), .C(_7294_), .Y(_7299_) );
NAND3X1 NAND3X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_7297_), .B(_7298_), .C(_7299_), .Y(_7300_) );
NAND3X1 NAND3X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_5267_), .B(_7296_), .C(_7300_), .Y(_7301_) );
AOI21X1 AOI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_7298_), .B(_7299_), .C(_7297_), .Y(_7302_) );
AOI21X1 AOI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_7290_), .B(_7295_), .C(_7134_), .Y(_7304_) );
OAI21X1 OAI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_7304_), .C(_5266_), .Y(_7305_) );
NAND3X1 NAND3X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_5613_), .B(_7301_), .C(_7305_), .Y(_7306_) );
NAND2X1 NAND2X1_923 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_158_), .B(_7306_), .Y(_7307_) );
INVX1 INVX1_949 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_158_), .Y(_7308_) );
NAND2X1 NAND2X1_924 ( .gnd(gnd), .vdd(vdd), .A(_7296_), .B(_7300_), .Y(_7309_) );
AOI21X1 AOI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_5266_), .B(_7309_), .C(_5614_), .Y(_7310_) );
NAND3X1 NAND3X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_7308_), .B(_7301_), .C(_7310_), .Y(_7311_) );
NAND3X1 NAND3X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_7133_), .B(_7311_), .C(_7307_), .Y(_7312_) );
NAND3X1 NAND3X1_1688 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_158_), .B(_7301_), .C(_7310_), .Y(_7313_) );
NAND2X1 NAND2X1_925 ( .gnd(gnd), .vdd(vdd), .A(_7308_), .B(_7306_), .Y(_7315_) );
NAND3X1 NAND3X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_6970_), .B(_7313_), .C(_7315_), .Y(_7316_) );
AOI21X1 AOI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_7312_), .B(_7316_), .C(_7132_), .Y(_7317_) );
NAND3X1 NAND3X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_6970_), .B(_7311_), .C(_7307_), .Y(_7318_) );
NAND3X1 NAND3X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_7133_), .B(_7313_), .C(_7315_), .Y(_7319_) );
AOI21X1 AOI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_7318_), .B(_7319_), .C(_7131_), .Y(_7320_) );
OAI21X1 OAI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .B(_7320_), .C(_7879_), .Y(_7321_) );
NAND3X1 NAND3X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_7131_), .B(_7318_), .C(_7319_), .Y(_7322_) );
NAND3X1 NAND3X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_7132_), .B(_7312_), .C(_7316_), .Y(_7323_) );
NAND3X1 NAND3X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_8092_), .B(_7322_), .C(_7323_), .Y(_7324_) );
NAND3X1 NAND3X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_5648_), .B(_7324_), .C(_7321_), .Y(_7326_) );
NAND2X1 NAND2X1_926 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_174_), .B(_7326_), .Y(_7327_) );
INVX1 INVX1_950 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_174_), .Y(_7328_) );
OAI21X1 OAI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .B(_7320_), .C(_8092_), .Y(_7329_) );
NAND3X1 NAND3X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_7879_), .B(_7322_), .C(_7323_), .Y(_7330_) );
NAND2X1 NAND2X1_927 ( .gnd(gnd), .vdd(vdd), .A(_7330_), .B(_7329_), .Y(_7331_) );
NAND3X1 NAND3X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_7328_), .B(_5648_), .C(_7331_), .Y(_7332_) );
NAND3X1 NAND3X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_7130_), .B(_7332_), .C(_7327_), .Y(_7333_) );
NAND3X1 NAND3X1_1699 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_174_), .B(_5648_), .C(_7331_), .Y(_7334_) );
NAND2X1 NAND2X1_928 ( .gnd(gnd), .vdd(vdd), .A(_7328_), .B(_7326_), .Y(_7335_) );
NAND3X1 NAND3X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_6992_), .B(_7334_), .C(_7335_), .Y(_7337_) );
AOI21X1 AOI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_7333_), .B(_7337_), .C(_7129_), .Y(_7338_) );
NAND3X1 NAND3X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_6992_), .B(_7332_), .C(_7327_), .Y(_7339_) );
NAND3X1 NAND3X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_7130_), .B(_7334_), .C(_7335_), .Y(_7340_) );
AOI21X1 AOI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_7339_), .B(_7340_), .C(_7128_), .Y(_7341_) );
OAI21X1 OAI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_7341_), .B(_7338_), .C(_7889_), .Y(_7342_) );
NAND3X1 NAND3X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_7128_), .B(_7339_), .C(_7340_), .Y(_7343_) );
NAND3X1 NAND3X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_7333_), .B(_7129_), .C(_7337_), .Y(_7344_) );
NAND3X1 NAND3X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_5261_), .B(_7343_), .C(_7344_), .Y(_7345_) );
NAND3X1 NAND3X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_5686_), .B(_7345_), .C(_7342_), .Y(_7346_) );
NAND2X1 NAND2X1_929 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_190_), .B(_7346_), .Y(_7348_) );
INVX1 INVX1_951 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_190_), .Y(_7349_) );
OAI21X1 OAI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_7341_), .B(_7338_), .C(_5261_), .Y(_7350_) );
NAND3X1 NAND3X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_7889_), .B(_7343_), .C(_7344_), .Y(_7351_) );
NAND2X1 NAND2X1_930 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .B(_7350_), .Y(_7352_) );
NAND3X1 NAND3X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_7349_), .B(_5686_), .C(_7352_), .Y(_7353_) );
NAND3X1 NAND3X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_7126_), .B(_7353_), .C(_7348_), .Y(_7354_) );
NAND3X1 NAND3X1_1710 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_190_), .B(_5686_), .C(_7352_), .Y(_7355_) );
NAND2X1 NAND2X1_931 ( .gnd(gnd), .vdd(vdd), .A(_7349_), .B(_7346_), .Y(_7356_) );
NAND3X1 NAND3X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_7022_), .B(_7355_), .C(_7356_), .Y(_7357_) );
AOI21X1 AOI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_7354_), .B(_7357_), .C(_7125_), .Y(_7359_) );
NAND3X1 NAND3X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_7022_), .B(_7353_), .C(_7348_), .Y(_7360_) );
NAND3X1 NAND3X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_7126_), .B(_7355_), .C(_7356_), .Y(_7361_) );
AOI21X1 AOI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_7360_), .B(_7361_), .C(_7124_), .Y(_7362_) );
OAI21X1 OAI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_7359_), .B(_7362_), .C(_5257_), .Y(_7363_) );
NAND3X1 NAND3X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(_7360_), .C(_7361_), .Y(_7364_) );
NAND3X1 NAND3X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_7354_), .B(_7357_), .C(_7125_), .Y(_7365_) );
NAND3X1 NAND3X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_5258_), .B(_7364_), .C(_7365_), .Y(_7366_) );
NAND3X1 NAND3X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_5722_), .B(_7366_), .C(_7363_), .Y(_7367_) );
NAND2X1 NAND2X1_932 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_206_), .B(_7367_), .Y(_7368_) );
INVX1 INVX1_952 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_206_), .Y(_7370_) );
NAND3X1 NAND3X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_5257_), .B(_7364_), .C(_7365_), .Y(_7371_) );
OAI21X1 OAI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_7359_), .B(_7362_), .C(_5258_), .Y(_7372_) );
NAND2X1 NAND2X1_933 ( .gnd(gnd), .vdd(vdd), .A(_7371_), .B(_7372_), .Y(_7373_) );
NAND3X1 NAND3X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_7370_), .B(_5722_), .C(_7373_), .Y(_7374_) );
NAND3X1 NAND3X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_7037_), .B(_7374_), .C(_7368_), .Y(_7375_) );
INVX1 INVX1_953 ( .gnd(gnd), .vdd(vdd), .A(_7037_), .Y(_7376_) );
NAND3X1 NAND3X1_1721 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_206_), .B(_5722_), .C(_7373_), .Y(_7377_) );
NAND2X1 NAND2X1_934 ( .gnd(gnd), .vdd(vdd), .A(_7370_), .B(_7367_), .Y(_7378_) );
NAND3X1 NAND3X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_7376_), .B(_7377_), .C(_7378_), .Y(_7379_) );
NAND3X1 NAND3X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_7123_), .B(_7375_), .C(_7379_), .Y(_7381_) );
AOI21X1 AOI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_7052_), .B(_7049_), .C(_7043_), .Y(_7382_) );
AOI21X1 AOI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_7377_), .B(_7378_), .C(_7376_), .Y(_7383_) );
AOI21X1 AOI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_7374_), .B(_7368_), .C(_7037_), .Y(_7384_) );
OAI21X1 OAI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_7383_), .B(_7384_), .C(_7382_), .Y(_7385_) );
NAND3X1 NAND3X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_5254_), .B(_7381_), .C(_7385_), .Y(_7386_) );
NOR3X1 NOR3X1_203 ( .gnd(gnd), .vdd(vdd), .A(_7383_), .B(_7382_), .C(_7384_), .Y(_7387_) );
AOI21X1 AOI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_7375_), .B(_7379_), .C(_7123_), .Y(_7388_) );
OAI21X1 OAI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_7387_), .B(_7388_), .C(_7907_), .Y(_7389_) );
NAND3X1 NAND3X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_5759_), .B(_7386_), .C(_7389_), .Y(_7390_) );
NAND2X1 NAND2X1_935 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_222_), .B(_7390_), .Y(_7392_) );
INVX1 INVX1_954 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_222_), .Y(_7393_) );
NAND2X1 NAND2X1_936 ( .gnd(gnd), .vdd(vdd), .A(_7381_), .B(_7385_), .Y(_7394_) );
AOI21X1 AOI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_7907_), .B(_7394_), .C(_5760_), .Y(_7395_) );
NAND3X1 NAND3X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_7393_), .B(_7386_), .C(_7395_), .Y(_7396_) );
NAND3X1 NAND3X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_7066_), .B(_7396_), .C(_7392_), .Y(_7397_) );
INVX1 INVX1_955 ( .gnd(gnd), .vdd(vdd), .A(_7066_), .Y(_7398_) );
NAND3X1 NAND3X1_1728 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_222_), .B(_7386_), .C(_7395_), .Y(_7399_) );
NAND2X1 NAND2X1_937 ( .gnd(gnd), .vdd(vdd), .A(_7393_), .B(_7390_), .Y(_7400_) );
NAND3X1 NAND3X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_7398_), .B(_7399_), .C(_7400_), .Y(_7401_) );
NAND3X1 NAND3X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_7122_), .B(_7397_), .C(_7401_), .Y(_7403_) );
AOI21X1 AOI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_7068_), .B(_6757_), .C(_7071_), .Y(_7404_) );
NAND3X1 NAND3X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_7398_), .B(_7396_), .C(_7392_), .Y(_7405_) );
NAND3X1 NAND3X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_7066_), .B(_7399_), .C(_7400_), .Y(_7406_) );
NAND3X1 NAND3X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_7404_), .B(_7405_), .C(_7406_), .Y(_7407_) );
NAND3X1 NAND3X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_5251_), .B(_7403_), .C(_7407_), .Y(_7408_) );
AOI21X1 AOI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_7405_), .B(_7406_), .C(_7404_), .Y(_7409_) );
AOI21X1 AOI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_7397_), .B(_7401_), .C(_7122_), .Y(_7410_) );
OAI21X1 OAI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_7409_), .B(_7410_), .C(_5250_), .Y(_7411_) );
NAND3X1 NAND3X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_5796_), .B(_7408_), .C(_7411_), .Y(_7412_) );
NAND2X1 NAND2X1_938 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_238_), .B(_7412_), .Y(_7414_) );
INVX1 INVX1_956 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_238_), .Y(_7415_) );
NAND2X1 NAND2X1_939 ( .gnd(gnd), .vdd(vdd), .A(_7403_), .B(_7407_), .Y(_7416_) );
AOI21X1 AOI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_5250_), .B(_7416_), .C(_5797_), .Y(_7417_) );
NAND3X1 NAND3X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_7415_), .B(_7408_), .C(_7417_), .Y(_7418_) );
NAND3X1 NAND3X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_7081_), .B(_7418_), .C(_7414_), .Y(_7419_) );
INVX2 INVX2_226 ( .gnd(gnd), .vdd(vdd), .A(_7081_), .Y(_7420_) );
NAND3X1 NAND3X1_1738 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_238_), .B(_7408_), .C(_7417_), .Y(_7421_) );
NAND2X1 NAND2X1_940 ( .gnd(gnd), .vdd(vdd), .A(_7415_), .B(_7412_), .Y(_7422_) );
NAND3X1 NAND3X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_7420_), .B(_7421_), .C(_7422_), .Y(_7423_) );
NAND3X1 NAND3X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_7419_), .B(_7423_), .C(_7121_), .Y(_7425_) );
AOI21X1 AOI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_7096_), .B(_7093_), .C(_7087_), .Y(_7426_) );
AOI21X1 AOI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_7421_), .B(_7422_), .C(_7420_), .Y(_7427_) );
AOI21X1 AOI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_7418_), .B(_7414_), .C(_7081_), .Y(_7428_) );
OAI21X1 OAI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_7427_), .B(_7428_), .C(_7426_), .Y(_7429_) );
NAND3X1 NAND3X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_8157_), .B(_7425_), .C(_7429_), .Y(_7430_) );
NAND3X1 NAND3X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_7420_), .B(_7418_), .C(_7414_), .Y(_7431_) );
NAND3X1 NAND3X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_7081_), .B(_7421_), .C(_7422_), .Y(_7432_) );
AOI21X1 AOI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_7431_), .B(_7432_), .C(_7426_), .Y(_7433_) );
AOI21X1 AOI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_7419_), .B(_7423_), .C(_7121_), .Y(_7434_) );
OAI21X1 OAI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_7433_), .B(_7434_), .C(_7929_), .Y(_7436_) );
NAND3X1 NAND3X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_5831_), .B(_7430_), .C(_7436_), .Y(_7437_) );
NAND2X1 NAND2X1_941 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_254_), .B(_7437_), .Y(_7438_) );
INVX1 INVX1_957 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_254_), .Y(_7439_) );
NAND2X1 NAND2X1_942 ( .gnd(gnd), .vdd(vdd), .A(_7425_), .B(_7429_), .Y(_7440_) );
AOI21X1 AOI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_7929_), .B(_7440_), .C(_5832_), .Y(_7441_) );
NAND3X1 NAND3X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_7439_), .B(_7430_), .C(_7441_), .Y(_7442_) );
NAND3X1 NAND3X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_7120_), .B(_7442_), .C(_7438_), .Y(_7443_) );
INVX1 INVX1_958 ( .gnd(gnd), .vdd(vdd), .A(_7443_), .Y(_7444_) );
AOI21X1 AOI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_7442_), .B(_7438_), .C(_7120_), .Y(_7445_) );
OAI21X1 OAI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_7444_), .B(_7445_), .C(_7119_), .Y(_7447_) );
INVX1 INVX1_959 ( .gnd(gnd), .vdd(vdd), .A(_7445_), .Y(_7448_) );
NAND3X1 NAND3X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .B(_7443_), .C(_7448_), .Y(_7449_) );
NAND2X1 NAND2X1_943 ( .gnd(gnd), .vdd(vdd), .A(_7447_), .B(_7449_), .Y(module_1_H_22_) );
OAI21X1 OAI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .B(_7445_), .C(_7443_), .Y(_7450_) );
AOI21X1 AOI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_7430_), .B(_7441_), .C(_7439_), .Y(_7451_) );
INVX1 INVX1_960 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_255_), .Y(_7452_) );
OAI21X1 OAI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_7426_), .B(_7428_), .C(_7419_), .Y(_7453_) );
INVX1 INVX1_961 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .Y(_7454_) );
NAND2X1 NAND2X1_944 ( .gnd(gnd), .vdd(vdd), .A(_7397_), .B(_7403_), .Y(_7455_) );
OAI21X1 OAI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_7384_), .B(_7382_), .C(_7375_), .Y(_7457_) );
NAND2X1 NAND2X1_945 ( .gnd(gnd), .vdd(vdd), .A(_7360_), .B(_7364_), .Y(_7458_) );
NAND2X1 NAND2X1_946 ( .gnd(gnd), .vdd(vdd), .A(_7339_), .B(_7343_), .Y(_7459_) );
INVX1 INVX1_962 ( .gnd(gnd), .vdd(vdd), .A(_7459_), .Y(_7460_) );
NAND2X1 NAND2X1_947 ( .gnd(gnd), .vdd(vdd), .A(_7318_), .B(_7322_), .Y(_7461_) );
NAND2X1 NAND2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_7290_), .B(_7296_), .Y(_7462_) );
NAND2X1 NAND2X1_949 ( .gnd(gnd), .vdd(vdd), .A(_7274_), .B(_7279_), .Y(_7463_) );
INVX1 INVX1_963 ( .gnd(gnd), .vdd(vdd), .A(_7463_), .Y(_7464_) );
INVX1 INVX1_964 ( .gnd(gnd), .vdd(vdd), .A(_7269_), .Y(_7465_) );
NOR2X1 NOR2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .B(_8065_), .Y(_7466_) );
NAND2X1 NAND2X1_950 ( .gnd(gnd), .vdd(vdd), .A(_7246_), .B(_7251_), .Y(_7468_) );
INVX1 INVX1_965 ( .gnd(gnd), .vdd(vdd), .A(_7468_), .Y(_7469_) );
OAI21X1 OAI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_7232_), .B(_7230_), .C(_7224_), .Y(_7470_) );
INVX1 INVX1_966 ( .gnd(gnd), .vdd(vdd), .A(_8045_), .Y(_7471_) );
NAND2X1 NAND2X1_951 ( .gnd(gnd), .vdd(vdd), .A(_7202_), .B(_7207_), .Y(_7472_) );
INVX1 INVX1_967 ( .gnd(gnd), .vdd(vdd), .A(_7472_), .Y(_7473_) );
NAND2X1 NAND2X1_952 ( .gnd(gnd), .vdd(vdd), .A(_7180_), .B(_7185_), .Y(_7474_) );
INVX1 INVX1_968 ( .gnd(gnd), .vdd(vdd), .A(_6083_), .Y(_7475_) );
XNOR2X1 XNOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_7175_), .B(_7475_), .Y(_7476_) );
INVX1 INVX1_969 ( .gnd(gnd), .vdd(vdd), .A(_7476_), .Y(_7477_) );
INVX1 INVX1_970 ( .gnd(gnd), .vdd(vdd), .A(_7142_), .Y(_7479_) );
NAND2X1 NAND2X1_953 ( .gnd(gnd), .vdd(vdd), .A(_7162_), .B(_7165_), .Y(_7480_) );
OAI21X1 OAI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_7480_), .B(_7479_), .C(_7162_), .Y(_7481_) );
INVX1 INVX1_971 ( .gnd(gnd), .vdd(vdd), .A(_7481_), .Y(_7482_) );
INVX1 INVX1_972 ( .gnd(gnd), .vdd(vdd), .A(_7157_), .Y(_7483_) );
OAI21X1 OAI21X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_6813_), .B(_6818_), .C(_7153_), .Y(_7484_) );
OAI21X1 OAI21X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_6807_), .B(_7152_), .C(_7484_), .Y(_7485_) );
INVX1 INVX1_973 ( .gnd(gnd), .vdd(vdd), .A(_7485_), .Y(_7486_) );
OAI21X1 OAI21X1_1169 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_12_), .B(module_1_W_13_), .C(module_1_W_14_), .Y(_7487_) );
XOR2X1 XOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_11_), .B(module_1_W_15_), .Y(_7488_) );
XNOR2X1 XNOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_7488_), .B(_7487_), .Y(_7490_) );
XOR2X1 XOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_7980_), .B(module_1_W_31_), .Y(_7491_) );
XNOR2X1 XNOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_7491_), .B(_7490_), .Y(_7492_) );
XOR2X1 XOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_7150_), .B(_7492_), .Y(_7493_) );
XNOR2X1 XNOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_7493_), .B(_5879_), .Y(_7494_) );
XNOR2X1 XNOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_6047_), .B(bloque_datos[15]), .Y(_7495_) );
XNOR2X1 XNOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_7494_), .B(_7495_), .Y(_7496_) );
NOR2X1 NOR2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_7486_), .B(_7496_), .Y(_7497_) );
NAND2X1 NAND2X1_954 ( .gnd(gnd), .vdd(vdd), .A(_7486_), .B(_7496_), .Y(_7498_) );
INVX1 INVX1_974 ( .gnd(gnd), .vdd(vdd), .A(_7498_), .Y(_7499_) );
OR2X2 OR2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_7499_), .B(_7497_), .Y(_7501_) );
NOR2X1 NOR2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_7483_), .B(_7501_), .Y(_7502_) );
INVX1 INVX1_975 ( .gnd(gnd), .vdd(vdd), .A(_7502_), .Y(_7503_) );
OAI21X1 OAI21X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_7499_), .B(_7497_), .C(_7483_), .Y(_7504_) );
XNOR2X1 XNOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_6061_), .B(_5885_), .Y(_7505_) );
INVX1 INVX1_976 ( .gnd(gnd), .vdd(vdd), .A(_7505_), .Y(_7506_) );
NAND3X1 NAND3X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_7504_), .B(_7506_), .C(_7503_), .Y(_7507_) );
AOI21X1 AOI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_7504_), .B(_7503_), .C(_7506_), .Y(_7508_) );
INVX1 INVX1_977 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .Y(_7509_) );
NAND2X1 NAND2X1_955 ( .gnd(gnd), .vdd(vdd), .A(_7507_), .B(_7509_), .Y(_7510_) );
NOR2X1 NOR2X1_506 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf3_), .B(_7510_), .Y(_7512_) );
AND2X2 AND2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_7510_), .B(bloque_datos_31_bF_buf2_), .Y(_7513_) );
NOR2X1 NOR2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_7512_), .B(_7513_), .Y(_7514_) );
NAND2X1 NAND2X1_956 ( .gnd(gnd), .vdd(vdd), .A(_7482_), .B(_7514_), .Y(_7515_) );
OAI21X1 OAI21X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_7513_), .B(_7512_), .C(_7481_), .Y(_7516_) );
XOR2X1 XOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_5900_), .B(bloque_datos_47_bF_buf3_), .Y(_7517_) );
NAND3X1 NAND3X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_7516_), .B(_7517_), .C(_7515_), .Y(_7518_) );
AND2X2 AND2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_7514_), .B(_7482_), .Y(_7519_) );
NOR2X1 NOR2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_7482_), .B(_7514_), .Y(_7520_) );
INVX1 INVX1_978 ( .gnd(gnd), .vdd(vdd), .A(_7517_), .Y(_7521_) );
OAI21X1 OAI21X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_7519_), .B(_7520_), .C(_7521_), .Y(_7523_) );
AOI21X1 AOI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_7518_), .B(_7523_), .C(_7477_), .Y(_7524_) );
INVX1 INVX1_979 ( .gnd(gnd), .vdd(vdd), .A(_7524_), .Y(_7525_) );
NAND3X1 NAND3X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_7477_), .B(_7518_), .C(_7523_), .Y(_7526_) );
NAND3X1 NAND3X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_7474_), .B(_7526_), .C(_7525_), .Y(_7527_) );
INVX1 INVX1_980 ( .gnd(gnd), .vdd(vdd), .A(_7474_), .Y(_7528_) );
INVX1 INVX1_981 ( .gnd(gnd), .vdd(vdd), .A(_7526_), .Y(_7529_) );
OAI21X1 OAI21X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_7529_), .B(_7524_), .C(_7528_), .Y(_7530_) );
OAI21X1 OAI21X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_5911_), .B(_5908_), .C(_8201_), .Y(_7531_) );
NAND2X1 NAND2X1_957 ( .gnd(gnd), .vdd(vdd), .A(_8030_), .B(_6035_), .Y(_7532_) );
NAND2X1 NAND2X1_958 ( .gnd(gnd), .vdd(vdd), .A(_7531_), .B(_7532_), .Y(_7534_) );
AOI21X1 AOI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_7530_), .B(_7527_), .C(_7534_), .Y(_7535_) );
NAND3X1 NAND3X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_7528_), .B(_7526_), .C(_7525_), .Y(_7536_) );
OAI21X1 OAI21X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_7529_), .B(_7524_), .C(_7474_), .Y(_7537_) );
AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_7531_), .B(_7532_), .C(_7536_), .D(_7537_), .Y(_7538_) );
NOR2X1 NOR2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_7535_), .B(_7538_), .Y(_7539_) );
XNOR2X1 XNOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_7197_), .B(bloque_datos[63]), .Y(_7540_) );
AND2X2 AND2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_7539_), .B(_7540_), .Y(_7541_) );
NOR2X1 NOR2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_7540_), .B(_7539_), .Y(_7542_) );
OAI21X1 OAI21X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_7541_), .B(_7542_), .C(_7473_), .Y(_7543_) );
NAND2X1 NAND2X1_959 ( .gnd(gnd), .vdd(vdd), .A(_7540_), .B(_7539_), .Y(_7545_) );
OR2X2 OR2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_7539_), .B(_7540_), .Y(_7546_) );
NAND3X1 NAND3X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_7472_), .B(_7545_), .C(_7546_), .Y(_7547_) );
NAND3X1 NAND3X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_7471_), .B(_7543_), .C(_7547_), .Y(_7548_) );
NAND3X1 NAND3X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_7473_), .B(_7545_), .C(_7546_), .Y(_7549_) );
OAI21X1 OAI21X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_7541_), .B(_7542_), .C(_7472_), .Y(_7550_) );
NAND3X1 NAND3X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_8045_), .B(_7550_), .C(_7549_), .Y(_7551_) );
NAND2X1 NAND2X1_960 ( .gnd(gnd), .vdd(vdd), .A(_7548_), .B(_7551_), .Y(_7552_) );
XOR2X1 XOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_6033_), .B(bloque_datos_79_bF_buf3_), .Y(_7553_) );
NOR2X1 NOR2X1_511 ( .gnd(gnd), .vdd(vdd), .A(_7219_), .B(_7553_), .Y(_7554_) );
INVX1 INVX1_982 ( .gnd(gnd), .vdd(vdd), .A(_7554_), .Y(_7556_) );
NAND2X1 NAND2X1_961 ( .gnd(gnd), .vdd(vdd), .A(_7219_), .B(_7553_), .Y(_7557_) );
NAND2X1 NAND2X1_962 ( .gnd(gnd), .vdd(vdd), .A(_7557_), .B(_7556_), .Y(_7558_) );
NAND2X1 NAND2X1_963 ( .gnd(gnd), .vdd(vdd), .A(_7558_), .B(_7552_), .Y(_7559_) );
OR2X2 OR2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_7552_), .B(_7558_), .Y(_7560_) );
NAND3X1 NAND3X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_7470_), .B(_7559_), .C(_7560_), .Y(_7561_) );
INVX1 INVX1_983 ( .gnd(gnd), .vdd(vdd), .A(_7470_), .Y(_7562_) );
AND2X2 AND2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_7552_), .B(_7558_), .Y(_7563_) );
NOR2X1 NOR2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_7558_), .B(_7552_), .Y(_7564_) );
OAI21X1 OAI21X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_7563_), .B(_7564_), .C(_7562_), .Y(_7565_) );
NOR2X1 NOR2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_8051_), .B(_8053_), .Y(_7567_) );
XNOR2X1 XNOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_6031_), .B(_7567_), .Y(_7568_) );
INVX1 INVX1_984 ( .gnd(gnd), .vdd(vdd), .A(_7568_), .Y(_7569_) );
AOI21X1 AOI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_7565_), .B(_7561_), .C(_7569_), .Y(_7570_) );
NAND3X1 NAND3X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_7562_), .B(_7559_), .C(_7560_), .Y(_7571_) );
OAI21X1 OAI21X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_7563_), .B(_7564_), .C(_7470_), .Y(_7572_) );
AOI21X1 AOI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_7572_), .B(_7571_), .C(_7568_), .Y(_7573_) );
NOR2X1 NOR2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_7570_), .B(_7573_), .Y(_7574_) );
NAND2X1 NAND2X1_964 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf3_), .B(_7241_), .Y(_7575_) );
NOR2X1 NOR2X1_515 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf2_), .B(_7241_), .Y(_7576_) );
INVX1 INVX1_985 ( .gnd(gnd), .vdd(vdd), .A(_7576_), .Y(_7578_) );
NAND2X1 NAND2X1_965 ( .gnd(gnd), .vdd(vdd), .A(_7575_), .B(_7578_), .Y(_7579_) );
NAND2X1 NAND2X1_966 ( .gnd(gnd), .vdd(vdd), .A(_7579_), .B(_7574_), .Y(_7580_) );
OR2X2 OR2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_7574_), .B(_7579_), .Y(_7581_) );
NAND3X1 NAND3X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_7469_), .B(_7580_), .C(_7581_), .Y(_7582_) );
AND2X2 AND2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_7574_), .B(_7579_), .Y(_7583_) );
NOR2X1 NOR2X1_516 ( .gnd(gnd), .vdd(vdd), .A(_7579_), .B(_7574_), .Y(_7584_) );
OAI21X1 OAI21X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_7583_), .B(_7584_), .C(_7468_), .Y(_7585_) );
AOI21X1 AOI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_7585_), .B(_7582_), .C(_7466_), .Y(_7586_) );
INVX1 INVX1_986 ( .gnd(gnd), .vdd(vdd), .A(_7466_), .Y(_7587_) );
OAI21X1 OAI21X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_7583_), .B(_7584_), .C(_7469_), .Y(_7589_) );
NAND3X1 NAND3X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_7468_), .B(_7580_), .C(_7581_), .Y(_7590_) );
AOI21X1 AOI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_7589_), .B(_7590_), .C(_7587_), .Y(_7591_) );
OAI21X1 OAI21X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_7586_), .B(_7591_), .C(_7465_), .Y(_7592_) );
NAND3X1 NAND3X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_7587_), .B(_7589_), .C(_7590_), .Y(_7593_) );
NAND3X1 NAND3X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_7466_), .B(_7585_), .C(_7582_), .Y(_7594_) );
NAND3X1 NAND3X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_7269_), .B(_7593_), .C(_7594_), .Y(_7595_) );
NAND2X1 NAND2X1_967 ( .gnd(gnd), .vdd(vdd), .A(_7595_), .B(_7592_), .Y(_7596_) );
AOI21X1 AOI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_7464_), .B(_7596_), .C(_5944_), .Y(_7597_) );
OAI21X1 OAI21X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_7464_), .B(_7596_), .C(_7597_), .Y(_7598_) );
XOR2X1 XOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_6200_), .B(module_1_W_143_), .Y(_7600_) );
XOR2X1 XOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_7598_), .B(_7600_), .Y(_7601_) );
XOR2X1 XOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_7601_), .B(_7284_), .Y(_7602_) );
NAND2X1 NAND2X1_968 ( .gnd(gnd), .vdd(vdd), .A(_7462_), .B(_7602_), .Y(_7603_) );
INVX1 INVX1_987 ( .gnd(gnd), .vdd(vdd), .A(_7462_), .Y(_7604_) );
XNOR2X1 XNOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_7601_), .B(_7284_), .Y(_7605_) );
AOI21X1 AOI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_7604_), .B(_7605_), .C(_6198_), .Y(_7606_) );
XNOR2X1 XNOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_8088_), .B(module_1_W_159_), .Y(_7607_) );
NAND3X1 NAND3X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_7603_), .B(_7607_), .C(_7606_), .Y(_7608_) );
NOR2X1 NOR2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_7604_), .B(_7605_), .Y(_7609_) );
OAI21X1 OAI21X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_7602_), .B(_7462_), .C(_5953_), .Y(_7611_) );
INVX1 INVX1_988 ( .gnd(gnd), .vdd(vdd), .A(_7607_), .Y(_7612_) );
OAI21X1 OAI21X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_7611_), .B(_7609_), .C(_7612_), .Y(_7613_) );
NAND2X1 NAND2X1_969 ( .gnd(gnd), .vdd(vdd), .A(_7608_), .B(_7613_), .Y(_7614_) );
XOR2X1 XOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_7614_), .B(_7307_), .Y(_7615_) );
NAND2X1 NAND2X1_970 ( .gnd(gnd), .vdd(vdd), .A(_7461_), .B(_7615_), .Y(_7616_) );
INVX1 INVX1_989 ( .gnd(gnd), .vdd(vdd), .A(_7461_), .Y(_7617_) );
XNOR2X1 XNOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_7614_), .B(_7307_), .Y(_7618_) );
AOI21X1 AOI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_7617_), .B(_7618_), .C(_5966_), .Y(_7619_) );
XOR2X1 XOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_8099_), .B(module_1_W_175_), .Y(_7620_) );
NAND3X1 NAND3X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_7616_), .B(_7620_), .C(_7619_), .Y(_7622_) );
NOR2X1 NOR2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_7617_), .B(_7618_), .Y(_7623_) );
OAI21X1 OAI21X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_7615_), .B(_7461_), .C(_6027_), .Y(_7624_) );
INVX1 INVX1_990 ( .gnd(gnd), .vdd(vdd), .A(_7620_), .Y(_7625_) );
OAI21X1 OAI21X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_7624_), .B(_7623_), .C(_7625_), .Y(_7626_) );
NAND2X1 NAND2X1_971 ( .gnd(gnd), .vdd(vdd), .A(_7622_), .B(_7626_), .Y(_7627_) );
XNOR2X1 XNOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_7627_), .B(_7327_), .Y(_7628_) );
NAND2X1 NAND2X1_972 ( .gnd(gnd), .vdd(vdd), .A(_7460_), .B(_7628_), .Y(_7629_) );
XOR2X1 XOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_7627_), .B(_7327_), .Y(_7630_) );
AOI21X1 AOI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_7459_), .B(_7630_), .C(_5976_), .Y(_7631_) );
AND2X2 AND2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_4681_), .B(module_1_W_191_), .Y(_7633_) );
NOR2X1 NOR2X1_519 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_191_), .B(_4681_), .Y(_7634_) );
NOR2X1 NOR2X1_520 ( .gnd(gnd), .vdd(vdd), .A(_7634_), .B(_7633_), .Y(_7635_) );
NAND3X1 NAND3X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_7629_), .B(_7635_), .C(_7631_), .Y(_7636_) );
NOR2X1 NOR2X1_521 ( .gnd(gnd), .vdd(vdd), .A(_7459_), .B(_7630_), .Y(_7637_) );
OAI21X1 OAI21X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_7628_), .B(_7460_), .C(_6023_), .Y(_7638_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_7633_), .B(_7634_), .C(_7638_), .D(_7637_), .Y(_7639_) );
NAND2X1 NAND2X1_973 ( .gnd(gnd), .vdd(vdd), .A(_7636_), .B(_7639_), .Y(_7640_) );
XOR2X1 XOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_7640_), .B(_7348_), .Y(_7641_) );
NAND2X1 NAND2X1_974 ( .gnd(gnd), .vdd(vdd), .A(_7458_), .B(_7641_), .Y(_7642_) );
INVX1 INVX1_991 ( .gnd(gnd), .vdd(vdd), .A(_7458_), .Y(_7644_) );
XNOR2X1 XNOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_7640_), .B(_7348_), .Y(_7645_) );
AOI21X1 AOI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_7644_), .B(_7645_), .C(_6262_), .Y(_7646_) );
OAI21X1 OAI21X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_8120_), .B(_8123_), .C(module_1_W_207_), .Y(_7647_) );
INVX1 INVX1_992 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_207_), .Y(_7648_) );
NAND3X1 NAND3X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_7648_), .B(_8122_), .C(_8127_), .Y(_7649_) );
NAND2X1 NAND2X1_975 ( .gnd(gnd), .vdd(vdd), .A(_7649_), .B(_7647_), .Y(_7650_) );
INVX1 INVX1_993 ( .gnd(gnd), .vdd(vdd), .A(_7650_), .Y(_7651_) );
NAND3X1 NAND3X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_7642_), .B(_7651_), .C(_7646_), .Y(_7652_) );
NOR2X1 NOR2X1_522 ( .gnd(gnd), .vdd(vdd), .A(_7644_), .B(_7645_), .Y(_7653_) );
OAI21X1 OAI21X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_7641_), .B(_7458_), .C(_5985_), .Y(_7655_) );
OAI21X1 OAI21X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_7655_), .B(_7653_), .C(_7650_), .Y(_7656_) );
NAND2X1 NAND2X1_976 ( .gnd(gnd), .vdd(vdd), .A(_7652_), .B(_7656_), .Y(_7657_) );
XOR2X1 XOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_7657_), .B(_7368_), .Y(_7658_) );
XNOR2X1 XNOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_7658_), .B(_7457_), .Y(_7659_) );
OAI21X1 OAI21X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_8135_), .B(_8138_), .C(module_1_W_223_), .Y(_7660_) );
INVX1 INVX1_994 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_223_), .Y(_7661_) );
NAND2X1 NAND2X1_977 ( .gnd(gnd), .vdd(vdd), .A(_7661_), .B(_8140_), .Y(_7662_) );
NAND2X1 NAND2X1_978 ( .gnd(gnd), .vdd(vdd), .A(_7660_), .B(_7662_), .Y(_7663_) );
NOR3X1 NOR3X1_204 ( .gnd(gnd), .vdd(vdd), .A(_7663_), .B(_5996_), .C(_7659_), .Y(_7664_) );
XOR2X1 XOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_7658_), .B(_7457_), .Y(_7666_) );
AND2X2 AND2X2_152 ( .gnd(gnd), .vdd(vdd), .A(_7662_), .B(_7660_), .Y(_7667_) );
AOI21X1 AOI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_6275_), .B(_7666_), .C(_7667_), .Y(_7668_) );
OAI21X1 OAI21X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_7664_), .B(_7668_), .C(_7392_), .Y(_7669_) );
INVX1 INVX1_995 ( .gnd(gnd), .vdd(vdd), .A(_7392_), .Y(_7670_) );
NAND3X1 NAND3X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_6275_), .B(_7666_), .C(_7667_), .Y(_7671_) );
OAI21X1 OAI21X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_7659_), .B(_5996_), .C(_7663_), .Y(_7672_) );
NAND3X1 NAND3X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_7670_), .B(_7671_), .C(_7672_), .Y(_7673_) );
AND2X2 AND2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_7669_), .B(_7673_), .Y(_7674_) );
NAND2X1 NAND2X1_979 ( .gnd(gnd), .vdd(vdd), .A(_7455_), .B(_7674_), .Y(_7675_) );
INVX1 INVX1_996 ( .gnd(gnd), .vdd(vdd), .A(_7455_), .Y(_7677_) );
NAND2X1 NAND2X1_980 ( .gnd(gnd), .vdd(vdd), .A(_7673_), .B(_7669_), .Y(_7678_) );
AOI21X1 AOI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_7678_), .B(_7677_), .C(_6006_), .Y(_7679_) );
OAI21X1 OAI21X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_8151_), .B(_8146_), .C(module_1_W_239_), .Y(_7680_) );
INVX1 INVX1_997 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_239_), .Y(_7681_) );
NAND3X1 NAND3X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_7681_), .B(_8145_), .C(_8150_), .Y(_7682_) );
AND2X2 AND2X2_154 ( .gnd(gnd), .vdd(vdd), .A(_7680_), .B(_7682_), .Y(_7683_) );
NAND3X1 NAND3X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_7675_), .B(_7679_), .C(_7683_), .Y(_7684_) );
NOR2X1 NOR2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_7678_), .B(_7677_), .Y(_7685_) );
OAI21X1 OAI21X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_7674_), .B(_7455_), .C(_6019_), .Y(_7686_) );
NAND2X1 NAND2X1_981 ( .gnd(gnd), .vdd(vdd), .A(_7682_), .B(_7680_), .Y(_7688_) );
OAI21X1 OAI21X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_7686_), .B(_7685_), .C(_7688_), .Y(_7689_) );
NAND2X1 NAND2X1_982 ( .gnd(gnd), .vdd(vdd), .A(_7689_), .B(_7684_), .Y(_7690_) );
XNOR2X1 XNOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_7690_), .B(_7414_), .Y(_7691_) );
NOR2X1 NOR2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_7454_), .B(_7691_), .Y(_7692_) );
XOR2X1 XOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_7690_), .B(_7414_), .Y(_7693_) );
OAI21X1 OAI21X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_7693_), .B(_7453_), .C(_6018_), .Y(_7694_) );
OAI21X1 OAI21X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_7694_), .B(_7692_), .C(_7452_), .Y(_7695_) );
OAI21X1 OAI21X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_7433_), .B(_7427_), .C(_7693_), .Y(_7696_) );
AOI21X1 AOI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_7454_), .B(_7691_), .C(_6017_), .Y(_7697_) );
NAND3X1 NAND3X1_1773 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_255_), .B(_7696_), .C(_7697_), .Y(_7699_) );
NAND3X1 NAND3X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_7451_), .B(_7699_), .C(_7695_), .Y(_7700_) );
NAND3X1 NAND3X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_7452_), .B(_7696_), .C(_7697_), .Y(_7701_) );
OAI21X1 OAI21X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_7694_), .B(_7692_), .C(module_1_W_255_), .Y(_7702_) );
NAND3X1 NAND3X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_7438_), .B(_7701_), .C(_7702_), .Y(_7703_) );
NAND2X1 NAND2X1_983 ( .gnd(gnd), .vdd(vdd), .A(_7703_), .B(_7700_), .Y(_7704_) );
XNOR2X1 XNOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_7450_), .B(_7704_), .Y(module_1_H_23_) );
INVX1 INVX1_998 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_241_), .Y(_6254_) );
AND2X2 AND2X2_155 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_0_), .B(module_1_W_16_), .Y(_6265_) );
NOR2X1 NOR2X1_525 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_0_), .B(module_1_W_16_), .Y(_6276_) );
OAI21X1 OAI21X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_6265_), .B(_6276_), .C(bloque_datos[0]), .Y(_6287_) );
INVX1 INVX1_999 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(_6298_) );
NOR2X1 NOR2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_6276_), .B(_6265_), .Y(_6309_) );
NAND2X1 NAND2X1_984 ( .gnd(gnd), .vdd(vdd), .A(_6298_), .B(_6309_), .Y(_6320_) );
NAND2X1 NAND2X1_985 ( .gnd(gnd), .vdd(vdd), .A(_6287_), .B(_6320_), .Y(_6331_) );
NAND2X1 NAND2X1_986 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf3_), .B(_6331_), .Y(_6342_) );
OR2X2 OR2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_6331_), .B(bloque_datos_16_bF_buf2_), .Y(_6353_) );
NAND2X1 NAND2X1_987 ( .gnd(gnd), .vdd(vdd), .A(_6342_), .B(_6353_), .Y(_6362_) );
NAND2X1 NAND2X1_988 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf3_), .B(_6362_), .Y(_6371_) );
OR2X2 OR2X2_152 ( .gnd(gnd), .vdd(vdd), .A(_6362_), .B(bloque_datos_32_bF_buf2_), .Y(_6381_) );
NAND2X1 NAND2X1_989 ( .gnd(gnd), .vdd(vdd), .A(_6371_), .B(_6381_), .Y(_6392_) );
NAND2X1 NAND2X1_990 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_48_bF_buf3_), .B(_6392_), .Y(_6403_) );
OR2X2 OR2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_6392_), .B(bloque_datos_48_bF_buf2_), .Y(_6414_) );
NAND2X1 NAND2X1_991 ( .gnd(gnd), .vdd(vdd), .A(_6403_), .B(_6414_), .Y(_6425_) );
NAND2X1 NAND2X1_992 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_64_bF_buf3_), .B(_6425_), .Y(_6436_) );
OR2X2 OR2X2_154 ( .gnd(gnd), .vdd(vdd), .A(_6425_), .B(bloque_datos_64_bF_buf2_), .Y(_6447_) );
NAND2X1 NAND2X1_993 ( .gnd(gnd), .vdd(vdd), .A(_6436_), .B(_6447_), .Y(_6458_) );
NAND2X1 NAND2X1_994 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf3_), .B(_6458_), .Y(_6469_) );
OR2X2 OR2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_6458_), .B(bloque_datos_80_bF_buf2_), .Y(_6480_) );
NAND2X1 NAND2X1_995 ( .gnd(gnd), .vdd(vdd), .A(_6469_), .B(_6480_), .Y(_6491_) );
NAND2X1 NAND2X1_996 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_128_), .B(_6491_), .Y(_6502_) );
OR2X2 OR2X2_156 ( .gnd(gnd), .vdd(vdd), .A(_6491_), .B(module_1_W_128_), .Y(_6513_) );
NAND2X1 NAND2X1_997 ( .gnd(gnd), .vdd(vdd), .A(_6502_), .B(_6513_), .Y(_6524_) );
NAND2X1 NAND2X1_998 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_144_), .B(_6524_), .Y(_6535_) );
OR2X2 OR2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_6524_), .B(module_1_W_144_), .Y(_6546_) );
NAND2X1 NAND2X1_999 ( .gnd(gnd), .vdd(vdd), .A(_6535_), .B(_6546_), .Y(_6557_) );
NAND2X1 NAND2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_160_), .B(_6557_), .Y(_6568_) );
OR2X2 OR2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_6557_), .B(module_1_W_160_), .Y(_6579_) );
NAND2X1 NAND2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_6568_), .B(_6579_), .Y(_6590_) );
NAND2X1 NAND2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_176_), .B(_6590_), .Y(_6601_) );
OR2X2 OR2X2_159 ( .gnd(gnd), .vdd(vdd), .A(_6590_), .B(module_1_W_176_), .Y(_6612_) );
NAND2X1 NAND2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_6601_), .B(_6612_), .Y(_6623_) );
NAND2X1 NAND2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_192_), .B(_6623_), .Y(_6634_) );
OR2X2 OR2X2_160 ( .gnd(gnd), .vdd(vdd), .A(_6623_), .B(module_1_W_192_), .Y(_6645_) );
NAND2X1 NAND2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_6634_), .B(_6645_), .Y(_6656_) );
NAND2X1 NAND2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_208_), .B(_6656_), .Y(_6667_) );
OR2X2 OR2X2_161 ( .gnd(gnd), .vdd(vdd), .A(_6656_), .B(module_1_W_208_), .Y(_6678_) );
NAND2X1 NAND2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_6667_), .B(_6678_), .Y(_6689_) );
INVX2 INVX2_227 ( .gnd(gnd), .vdd(vdd), .A(_6689_), .Y(_6700_) );
NOR2X1 NOR2X1_527 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_224_), .B(_6700_), .Y(_6711_) );
INVX1 INVX1_1000 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_225_), .Y(_6722_) );
INVX2 INVX2_228 ( .gnd(gnd), .vdd(vdd), .A(_6656_), .Y(_6733_) );
NOR2X1 NOR2X1_528 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_208_), .B(_6733_), .Y(_6744_) );
INVX2 INVX2_229 ( .gnd(gnd), .vdd(vdd), .A(_6623_), .Y(_6754_) );
NOR2X1 NOR2X1_529 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_192_), .B(_6754_), .Y(_6765_) );
INVX1 INVX1_1001 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_193_), .Y(_6776_) );
INVX2 INVX2_230 ( .gnd(gnd), .vdd(vdd), .A(_6590_), .Y(_6787_) );
NOR2X1 NOR2X1_530 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_176_), .B(_6787_), .Y(_6798_) );
INVX2 INVX2_231 ( .gnd(gnd), .vdd(vdd), .A(_6557_), .Y(_6809_) );
NOR2X1 NOR2X1_531 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_160_), .B(_6809_), .Y(_6820_) );
INVX1 INVX1_1002 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_161_), .Y(_6831_) );
INVX2 INVX2_232 ( .gnd(gnd), .vdd(vdd), .A(_6524_), .Y(_6842_) );
NOR2X1 NOR2X1_532 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_144_), .B(_6842_), .Y(_6853_) );
INVX1 INVX1_1003 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_145_), .Y(_6864_) );
INVX2 INVX2_233 ( .gnd(gnd), .vdd(vdd), .A(_6491_), .Y(_6875_) );
NOR2X1 NOR2X1_533 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_128_), .B(_6875_), .Y(_6886_) );
INVX2 INVX2_234 ( .gnd(gnd), .vdd(vdd), .A(_6458_), .Y(_6897_) );
NOR2X1 NOR2X1_534 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf1_), .B(_6897_), .Y(_6908_) );
AOI21X1 AOI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_6403_), .B(_6414_), .C(bloque_datos_64_bF_buf1_), .Y(_6919_) );
AOI21X1 AOI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_6371_), .B(_6381_), .C(bloque_datos_48_bF_buf1_), .Y(_6930_) );
INVX1 INVX1_1004 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_49_bF_buf3_), .Y(_6941_) );
AOI21X1 AOI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_6342_), .B(_6353_), .C(bloque_datos_32_bF_buf1_), .Y(_6952_) );
INVX1 INVX1_1005 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf2_), .Y(_6963_) );
AOI21X1 AOI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_6287_), .B(_6320_), .C(bloque_datos_16_bF_buf1_), .Y(_6974_) );
OAI21X1 OAI21X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_6265_), .B(_6276_), .C(_6298_), .Y(_6985_) );
INVX1 INVX1_1006 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(_6996_) );
INVX2 INVX2_235 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_0_), .Y(_7007_) );
NOR2X1 NOR2X1_535 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_16_), .B(_7007_), .Y(_7018_) );
NAND2X1 NAND2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_0_), .B(module_1_W_1_), .Y(_7029_) );
OR2X2 OR2X2_162 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_0_), .B(module_1_W_1_), .Y(_7040_) );
AOI21X1 AOI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_7029_), .B(_7040_), .C(module_1_W_17_), .Y(_7051_) );
INVX1 INVX1_1007 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_17_), .Y(_7062_) );
AND2X2 AND2X2_156 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_0_), .B(module_1_W_1_), .Y(_7073_) );
NOR2X1 NOR2X1_536 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_0_), .B(module_1_W_1_), .Y(_7084_) );
NOR3X1 NOR3X1_205 ( .gnd(gnd), .vdd(vdd), .A(_7062_), .B(_7084_), .C(_7073_), .Y(_7095_) );
OAI21X1 OAI21X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_7095_), .B(_7051_), .C(_7018_), .Y(_7106_) );
INVX1 INVX1_1008 ( .gnd(gnd), .vdd(vdd), .A(_7018_), .Y(_7116_) );
OAI21X1 OAI21X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_7073_), .B(_7084_), .C(_7062_), .Y(_7127_) );
NAND3X1 NAND3X1_1777 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_17_), .B(_7029_), .C(_7040_), .Y(_7138_) );
NAND3X1 NAND3X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_7127_), .B(_7138_), .C(_7116_), .Y(_7149_) );
NAND2X1 NAND2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_7149_), .B(_7106_), .Y(_7160_) );
NAND2X1 NAND2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_6996_), .B(_7160_), .Y(_7171_) );
OR2X2 OR2X2_163 ( .gnd(gnd), .vdd(vdd), .A(_7160_), .B(_6996_), .Y(_7182_) );
NAND2X1 NAND2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_7171_), .B(_7182_), .Y(_7193_) );
XNOR2X1 XNOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_7193_), .B(_6985_), .Y(_7204_) );
XNOR2X1 XNOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_7204_), .B(bloque_datos[17]), .Y(_7215_) );
AND2X2 AND2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_7215_), .B(_6974_), .Y(_7226_) );
NOR2X1 NOR2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_6974_), .B(_7215_), .Y(_7237_) );
OAI21X1 OAI21X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_7226_), .B(_7237_), .C(_6963_), .Y(_7248_) );
OR2X2 OR2X2_164 ( .gnd(gnd), .vdd(vdd), .A(_7226_), .B(_7237_), .Y(_7259_) );
NOR2X1 NOR2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_6963_), .B(_7259_), .Y(_7270_) );
INVX1 INVX1_1009 ( .gnd(gnd), .vdd(vdd), .A(_7270_), .Y(_7281_) );
NAND2X1 NAND2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_7248_), .B(_7281_), .Y(_7292_) );
AND2X2 AND2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_7292_), .B(_6952_), .Y(_7303_) );
NOR2X1 NOR2X1_539 ( .gnd(gnd), .vdd(vdd), .A(_6952_), .B(_7292_), .Y(_7314_) );
OAI21X1 OAI21X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(_7314_), .C(_6941_), .Y(_7325_) );
OR2X2 OR2X2_165 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(_7314_), .Y(_7336_) );
NOR2X1 NOR2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_6941_), .B(_7336_), .Y(_7347_) );
INVX1 INVX1_1010 ( .gnd(gnd), .vdd(vdd), .A(_7347_), .Y(_7358_) );
NAND2X1 NAND2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_7325_), .B(_7358_), .Y(_7369_) );
AND2X2 AND2X2_159 ( .gnd(gnd), .vdd(vdd), .A(_7369_), .B(_6930_), .Y(_7380_) );
NOR2X1 NOR2X1_541 ( .gnd(gnd), .vdd(vdd), .A(_6930_), .B(_7369_), .Y(_7391_) );
NOR2X1 NOR2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_7391_), .B(_7380_), .Y(_7402_) );
XNOR2X1 XNOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_7402_), .B(bloque_datos_65_bF_buf2_), .Y(_7413_) );
AND2X2 AND2X2_160 ( .gnd(gnd), .vdd(vdd), .A(_7413_), .B(_6919_), .Y(_7424_) );
NOR2X1 NOR2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_6919_), .B(_7413_), .Y(_7435_) );
NOR2X1 NOR2X1_544 ( .gnd(gnd), .vdd(vdd), .A(_7435_), .B(_7424_), .Y(_7446_) );
NOR2X1 NOR2X1_545 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf3_), .B(_7446_), .Y(_7456_) );
INVX1 INVX1_1011 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf2_), .Y(_7467_) );
INVX1 INVX1_1012 ( .gnd(gnd), .vdd(vdd), .A(_7446_), .Y(_7478_) );
NOR2X1 NOR2X1_546 ( .gnd(gnd), .vdd(vdd), .A(_7467_), .B(_7478_), .Y(_7489_) );
OAI21X1 OAI21X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_7489_), .B(_7456_), .C(_6908_), .Y(_7500_) );
OR2X2 OR2X2_166 ( .gnd(gnd), .vdd(vdd), .A(_7489_), .B(_7456_), .Y(_7511_) );
NOR2X1 NOR2X1_547 ( .gnd(gnd), .vdd(vdd), .A(_6908_), .B(_7511_), .Y(_7522_) );
INVX2 INVX2_236 ( .gnd(gnd), .vdd(vdd), .A(_7522_), .Y(_7533_) );
NAND2X1 NAND2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_7500_), .B(_7533_), .Y(_7544_) );
INVX2 INVX2_237 ( .gnd(gnd), .vdd(vdd), .A(_7544_), .Y(_7555_) );
NOR2X1 NOR2X1_548 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_129_), .B(_7555_), .Y(_7566_) );
AND2X2 AND2X2_161 ( .gnd(gnd), .vdd(vdd), .A(_7555_), .B(module_1_W_129_), .Y(_7577_) );
OAI21X1 OAI21X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_7577_), .B(_7566_), .C(_6886_), .Y(_7588_) );
OR2X2 OR2X2_167 ( .gnd(gnd), .vdd(vdd), .A(_7577_), .B(_7566_), .Y(_7599_) );
OR2X2 OR2X2_168 ( .gnd(gnd), .vdd(vdd), .A(_7599_), .B(_6886_), .Y(_7610_) );
NAND2X1 NAND2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_7588_), .B(_7610_), .Y(_7621_) );
NAND2X1 NAND2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_6864_), .B(_7621_), .Y(_7632_) );
NOR2X1 NOR2X1_549 ( .gnd(gnd), .vdd(vdd), .A(_6864_), .B(_7621_), .Y(_7643_) );
INVX1 INVX1_1013 ( .gnd(gnd), .vdd(vdd), .A(_7643_), .Y(_7654_) );
NAND2X1 NAND2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_7632_), .B(_7654_), .Y(_7665_) );
NAND2X1 NAND2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_6853_), .B(_7665_), .Y(_7676_) );
NOR2X1 NOR2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_6853_), .B(_7665_), .Y(_7687_) );
INVX1 INVX1_1014 ( .gnd(gnd), .vdd(vdd), .A(_7687_), .Y(_7698_) );
NAND2X1 NAND2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_7676_), .B(_7698_), .Y(_7705_) );
NAND2X1 NAND2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_6831_), .B(_7705_), .Y(_7706_) );
NOR2X1 NOR2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_6831_), .B(_7705_), .Y(_7707_) );
INVX1 INVX1_1015 ( .gnd(gnd), .vdd(vdd), .A(_7707_), .Y(_7708_) );
NAND2X1 NAND2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_7706_), .B(_7708_), .Y(_7709_) );
NAND2X1 NAND2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_6820_), .B(_7709_), .Y(_7710_) );
NOR2X1 NOR2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_6820_), .B(_7709_), .Y(_7711_) );
INVX1 INVX1_1016 ( .gnd(gnd), .vdd(vdd), .A(_7711_), .Y(_7712_) );
NAND2X1 NAND2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_7710_), .B(_7712_), .Y(_7713_) );
INVX2 INVX2_238 ( .gnd(gnd), .vdd(vdd), .A(_7713_), .Y(_7714_) );
NOR2X1 NOR2X1_553 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_177_), .B(_7714_), .Y(_7715_) );
NAND2X1 NAND2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_177_), .B(_7714_), .Y(_7716_) );
INVX2 INVX2_239 ( .gnd(gnd), .vdd(vdd), .A(_7716_), .Y(_7717_) );
OAI21X1 OAI21X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_7717_), .B(_7715_), .C(_6798_), .Y(_7718_) );
OR2X2 OR2X2_169 ( .gnd(gnd), .vdd(vdd), .A(_7717_), .B(_7715_), .Y(_7719_) );
NOR2X1 NOR2X1_554 ( .gnd(gnd), .vdd(vdd), .A(_6798_), .B(_7719_), .Y(_7720_) );
INVX1 INVX1_1017 ( .gnd(gnd), .vdd(vdd), .A(_7720_), .Y(_7721_) );
NAND2X1 NAND2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_7718_), .B(_7721_), .Y(_7722_) );
NAND2X1 NAND2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_6776_), .B(_7722_), .Y(_7723_) );
NOR2X1 NOR2X1_555 ( .gnd(gnd), .vdd(vdd), .A(_6776_), .B(_7722_), .Y(_7724_) );
INVX1 INVX1_1018 ( .gnd(gnd), .vdd(vdd), .A(_7724_), .Y(_7725_) );
NAND2X1 NAND2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_7723_), .B(_7725_), .Y(_7726_) );
NAND2X1 NAND2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_6765_), .B(_7726_), .Y(_7727_) );
NOR2X1 NOR2X1_556 ( .gnd(gnd), .vdd(vdd), .A(_6765_), .B(_7726_), .Y(_7728_) );
INVX1 INVX1_1019 ( .gnd(gnd), .vdd(vdd), .A(_7728_), .Y(_7729_) );
NAND2X1 NAND2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_7727_), .B(_7729_), .Y(_7730_) );
INVX2 INVX2_240 ( .gnd(gnd), .vdd(vdd), .A(_7730_), .Y(_7731_) );
NOR2X1 NOR2X1_557 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_209_), .B(_7731_), .Y(_7732_) );
NAND2X1 NAND2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_209_), .B(_7731_), .Y(_7733_) );
INVX2 INVX2_241 ( .gnd(gnd), .vdd(vdd), .A(_7733_), .Y(_7734_) );
OAI21X1 OAI21X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_7734_), .B(_7732_), .C(_6744_), .Y(_7735_) );
OR2X2 OR2X2_170 ( .gnd(gnd), .vdd(vdd), .A(_7734_), .B(_7732_), .Y(_7736_) );
NOR2X1 NOR2X1_558 ( .gnd(gnd), .vdd(vdd), .A(_6744_), .B(_7736_), .Y(_7737_) );
INVX2 INVX2_242 ( .gnd(gnd), .vdd(vdd), .A(_7737_), .Y(_7738_) );
NAND2X1 NAND2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_7735_), .B(_7738_), .Y(_7739_) );
NAND2X1 NAND2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_6722_), .B(_7739_), .Y(_7740_) );
NOR2X1 NOR2X1_559 ( .gnd(gnd), .vdd(vdd), .A(_6722_), .B(_7739_), .Y(_7741_) );
INVX1 INVX1_1020 ( .gnd(gnd), .vdd(vdd), .A(_7741_), .Y(_7742_) );
NAND2X1 NAND2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_7740_), .B(_7742_), .Y(_7743_) );
NAND2X1 NAND2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_6711_), .B(_7743_), .Y(_7744_) );
NOR2X1 NOR2X1_560 ( .gnd(gnd), .vdd(vdd), .A(_6711_), .B(_7743_), .Y(_7745_) );
INVX1 INVX1_1021 ( .gnd(gnd), .vdd(vdd), .A(_7745_), .Y(_7746_) );
NAND2X1 NAND2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_7744_), .B(_7746_), .Y(_7747_) );
NOR2X1 NOR2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_6254_), .B(_7747_), .Y(_7748_) );
INVX1 INVX1_1022 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_242_), .Y(_7749_) );
INVX1 INVX1_1023 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_194_), .Y(_7750_) );
INVX1 INVX1_1024 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_178_), .Y(_7751_) );
INVX1 INVX1_1025 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_162_), .Y(_7752_) );
NOR2X1 NOR2X1_562 ( .gnd(gnd), .vdd(vdd), .A(_6886_), .B(_7599_), .Y(_7753_) );
AND2X2 AND2X2_162 ( .gnd(gnd), .vdd(vdd), .A(_7402_), .B(bloque_datos_65_bF_buf1_), .Y(_7754_) );
INVX1 INVX1_1026 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf3_), .Y(_7755_) );
INVX1 INVX1_1027 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf3_), .Y(_7756_) );
INVX1 INVX1_1028 ( .gnd(gnd), .vdd(vdd), .A(_7237_), .Y(_7757_) );
NAND2X1 NAND2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .B(_7204_), .Y(_7758_) );
INVX1 INVX1_1029 ( .gnd(gnd), .vdd(vdd), .A(_6985_), .Y(_7759_) );
NOR2X1 NOR2X1_563 ( .gnd(gnd), .vdd(vdd), .A(_7759_), .B(_7193_), .Y(_7760_) );
INVX1 INVX1_1030 ( .gnd(gnd), .vdd(vdd), .A(_7182_), .Y(_7761_) );
INVX1 INVX1_1031 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf3_), .Y(_7762_) );
INVX1 INVX1_1032 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_18_), .Y(_7763_) );
NAND3X1 NAND3X1_1779 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_2_), .B(module_1_W_0_), .C(module_1_W_1_), .Y(_7764_) );
INVX2 INVX2_243 ( .gnd(gnd), .vdd(vdd), .A(_7764_), .Y(_7765_) );
AOI21X1 AOI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_0_), .B(module_1_W_1_), .C(module_1_W_2_), .Y(_7766_) );
OAI21X1 OAI21X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_7765_), .B(_7766_), .C(_7763_), .Y(_7767_) );
INVX2 INVX2_244 ( .gnd(gnd), .vdd(vdd), .A(_7766_), .Y(_7768_) );
NAND3X1 NAND3X1_1780 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_18_), .B(_7764_), .C(_7768_), .Y(_7769_) );
NAND3X1 NAND3X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_7095_), .B(_7769_), .C(_7767_), .Y(_7770_) );
AOI21X1 AOI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_7764_), .B(_7768_), .C(module_1_W_18_), .Y(_7771_) );
NOR3X1 NOR3X1_206 ( .gnd(gnd), .vdd(vdd), .A(_7763_), .B(_7766_), .C(_7765_), .Y(_7772_) );
OAI21X1 OAI21X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_7772_), .B(_7771_), .C(_7138_), .Y(_7773_) );
NAND2X1 NAND2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_7770_), .B(_7773_), .Y(_7774_) );
NOR2X1 NOR2X1_564 ( .gnd(gnd), .vdd(vdd), .A(_7149_), .B(_7774_), .Y(_7775_) );
INVX1 INVX1_1033 ( .gnd(gnd), .vdd(vdd), .A(_7149_), .Y(_7776_) );
AOI21X1 AOI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_7770_), .B(_7773_), .C(_7776_), .Y(_7777_) );
OAI21X1 OAI21X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_7775_), .B(_7777_), .C(_7762_), .Y(_7778_) );
OR2X2 OR2X2_171 ( .gnd(gnd), .vdd(vdd), .A(_7774_), .B(_7149_), .Y(_7779_) );
INVX1 INVX1_1034 ( .gnd(gnd), .vdd(vdd), .A(_7777_), .Y(_7780_) );
NAND3X1 NAND3X1_1782 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf2_), .B(_7780_), .C(_7779_), .Y(_7781_) );
NAND3X1 NAND3X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_7761_), .B(_7778_), .C(_7781_), .Y(_7782_) );
AOI21X1 AOI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_7780_), .B(_7779_), .C(bloque_datos_2_bF_buf1_), .Y(_7783_) );
NOR3X1 NOR3X1_207 ( .gnd(gnd), .vdd(vdd), .A(_7762_), .B(_7777_), .C(_7775_), .Y(_7784_) );
OAI21X1 OAI21X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_7783_), .B(_7784_), .C(_7182_), .Y(_7785_) );
NAND3X1 NAND3X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_7760_), .B(_7782_), .C(_7785_), .Y(_7786_) );
AOI21X1 AOI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_7782_), .B(_7785_), .C(_7760_), .Y(_7787_) );
INVX1 INVX1_1035 ( .gnd(gnd), .vdd(vdd), .A(_7787_), .Y(_7788_) );
AOI21X1 AOI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_7786_), .B(_7788_), .C(bloque_datos[18]), .Y(_7789_) );
INVX1 INVX1_1036 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .Y(_7790_) );
INVX1 INVX1_1037 ( .gnd(gnd), .vdd(vdd), .A(_7760_), .Y(_7791_) );
NOR3X1 NOR3X1_208 ( .gnd(gnd), .vdd(vdd), .A(_7784_), .B(_7182_), .C(_7783_), .Y(_7792_) );
AOI21X1 AOI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_7778_), .B(_7781_), .C(_7761_), .Y(_7793_) );
NOR3X1 NOR3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_7791_), .B(_7793_), .C(_7792_), .Y(_7794_) );
NOR3X1 NOR3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_7790_), .B(_7787_), .C(_7794_), .Y(_7795_) );
NOR3X1 NOR3X1_211 ( .gnd(gnd), .vdd(vdd), .A(_7758_), .B(_7795_), .C(_7789_), .Y(_7796_) );
INVX1 INVX1_1038 ( .gnd(gnd), .vdd(vdd), .A(_7758_), .Y(_7797_) );
OAI21X1 OAI21X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_7794_), .B(_7787_), .C(_7790_), .Y(_7798_) );
INVX2 INVX2_245 ( .gnd(gnd), .vdd(vdd), .A(_7795_), .Y(_7799_) );
AOI21X1 AOI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_7798_), .B(_7799_), .C(_7797_), .Y(_7800_) );
NOR3X1 NOR3X1_212 ( .gnd(gnd), .vdd(vdd), .A(_7757_), .B(_7796_), .C(_7800_), .Y(_7801_) );
NAND3X1 NAND3X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_7797_), .B(_7798_), .C(_7799_), .Y(_7802_) );
OAI21X1 OAI21X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_7789_), .B(_7795_), .C(_7758_), .Y(_7803_) );
AOI21X1 AOI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_7803_), .B(_7802_), .C(_7237_), .Y(_7804_) );
OAI21X1 OAI21X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_7801_), .B(_7804_), .C(_7756_), .Y(_7805_) );
NAND3X1 NAND3X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_7237_), .B(_7803_), .C(_7802_), .Y(_7806_) );
OAI21X1 OAI21X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_7800_), .B(_7796_), .C(_7757_), .Y(_7807_) );
NAND3X1 NAND3X1_1787 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf2_), .B(_7806_), .C(_7807_), .Y(_7808_) );
NAND3X1 NAND3X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_7270_), .B(_7808_), .C(_7805_), .Y(_7809_) );
AOI21X1 AOI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_7806_), .B(_7807_), .C(bloque_datos_34_bF_buf1_), .Y(_7810_) );
NOR3X1 NOR3X1_213 ( .gnd(gnd), .vdd(vdd), .A(_7756_), .B(_7804_), .C(_7801_), .Y(_7811_) );
OAI21X1 OAI21X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_7811_), .B(_7810_), .C(_7281_), .Y(_7812_) );
NAND3X1 NAND3X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_7314_), .B(_7809_), .C(_7812_), .Y(_7813_) );
AOI21X1 AOI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_7809_), .B(_7812_), .C(_7314_), .Y(_7814_) );
INVX1 INVX1_1039 ( .gnd(gnd), .vdd(vdd), .A(_7814_), .Y(_7815_) );
AOI21X1 AOI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_7813_), .B(_7815_), .C(bloque_datos_50_bF_buf2_), .Y(_7816_) );
INVX1 INVX1_1040 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_50_bF_buf1_), .Y(_7817_) );
INVX1 INVX1_1041 ( .gnd(gnd), .vdd(vdd), .A(_7813_), .Y(_7818_) );
NOR3X1 NOR3X1_214 ( .gnd(gnd), .vdd(vdd), .A(_7817_), .B(_7814_), .C(_7818_), .Y(_7819_) );
NOR2X1 NOR2X1_565 ( .gnd(gnd), .vdd(vdd), .A(_7816_), .B(_7819_), .Y(_7820_) );
NAND2X1 NAND2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_7347_), .B(_7820_), .Y(_7821_) );
OAI21X1 OAI21X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_7819_), .B(_7816_), .C(_7358_), .Y(_7822_) );
NAND3X1 NAND3X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_7391_), .B(_7822_), .C(_7821_), .Y(_7823_) );
INVX2 INVX2_246 ( .gnd(gnd), .vdd(vdd), .A(_7823_), .Y(_7824_) );
AOI21X1 AOI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_7822_), .B(_7821_), .C(_7391_), .Y(_7825_) );
OAI21X1 OAI21X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_7824_), .B(_7825_), .C(_7755_), .Y(_7826_) );
INVX1 INVX1_1042 ( .gnd(gnd), .vdd(vdd), .A(_7391_), .Y(_7827_) );
AND2X2 AND2X2_163 ( .gnd(gnd), .vdd(vdd), .A(_7820_), .B(_7347_), .Y(_7828_) );
INVX1 INVX1_1043 ( .gnd(gnd), .vdd(vdd), .A(_7822_), .Y(_7829_) );
OAI21X1 OAI21X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_7828_), .B(_7829_), .C(_7827_), .Y(_7830_) );
NAND3X1 NAND3X1_1791 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf2_), .B(_7823_), .C(_7830_), .Y(_7831_) );
NAND3X1 NAND3X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_7754_), .B(_7831_), .C(_7826_), .Y(_7832_) );
INVX1 INVX1_1044 ( .gnd(gnd), .vdd(vdd), .A(_7754_), .Y(_7833_) );
AOI21X1 AOI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_7823_), .B(_7830_), .C(bloque_datos_66_bF_buf1_), .Y(_7834_) );
NOR3X1 NOR3X1_215 ( .gnd(gnd), .vdd(vdd), .A(_7755_), .B(_7825_), .C(_7824_), .Y(_7835_) );
OAI21X1 OAI21X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_7835_), .B(_7834_), .C(_7833_), .Y(_7836_) );
NAND3X1 NAND3X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_7435_), .B(_7832_), .C(_7836_), .Y(_7837_) );
INVX2 INVX2_247 ( .gnd(gnd), .vdd(vdd), .A(_7435_), .Y(_7838_) );
NOR3X1 NOR3X1_216 ( .gnd(gnd), .vdd(vdd), .A(_7833_), .B(_7834_), .C(_7835_), .Y(_7839_) );
AOI21X1 AOI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_7831_), .B(_7826_), .C(_7754_), .Y(_7840_) );
OAI21X1 OAI21X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_7839_), .B(_7840_), .C(_7838_), .Y(_7841_) );
AOI21X1 AOI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_7837_), .B(_7841_), .C(bloque_datos_82_bF_buf2_), .Y(_7842_) );
INVX1 INVX1_1045 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf1_), .Y(_7843_) );
NOR3X1 NOR3X1_217 ( .gnd(gnd), .vdd(vdd), .A(_7838_), .B(_7840_), .C(_7839_), .Y(_7844_) );
AOI21X1 AOI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_7832_), .B(_7836_), .C(_7435_), .Y(_7845_) );
NOR3X1 NOR3X1_218 ( .gnd(gnd), .vdd(vdd), .A(_7843_), .B(_7845_), .C(_7844_), .Y(_7846_) );
NOR2X1 NOR2X1_566 ( .gnd(gnd), .vdd(vdd), .A(_7842_), .B(_7846_), .Y(_7847_) );
NAND2X1 NAND2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_7489_), .B(_7847_), .Y(_7848_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_7467_), .B(_7478_), .C(_7846_), .D(_7842_), .Y(_7849_) );
NAND3X1 NAND3X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_7522_), .B(_7849_), .C(_7848_), .Y(_7850_) );
AND2X2 AND2X2_164 ( .gnd(gnd), .vdd(vdd), .A(_7847_), .B(_7489_), .Y(_7851_) );
INVX2 INVX2_248 ( .gnd(gnd), .vdd(vdd), .A(_7849_), .Y(_7852_) );
OAI21X1 OAI21X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_7851_), .B(_7852_), .C(_7533_), .Y(_7853_) );
AOI21X1 AOI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_7850_), .B(_7853_), .C(module_1_W_130_), .Y(_7854_) );
INVX1 INVX1_1046 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_130_), .Y(_7855_) );
NOR3X1 NOR3X1_219 ( .gnd(gnd), .vdd(vdd), .A(_7852_), .B(_7533_), .C(_7851_), .Y(_7856_) );
AOI21X1 AOI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_7849_), .B(_7848_), .C(_7522_), .Y(_7857_) );
NOR3X1 NOR3X1_220 ( .gnd(gnd), .vdd(vdd), .A(_7855_), .B(_7857_), .C(_7856_), .Y(_7858_) );
NOR2X1 NOR2X1_567 ( .gnd(gnd), .vdd(vdd), .A(_7854_), .B(_7858_), .Y(_7859_) );
NAND2X1 NAND2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_7577_), .B(_7859_), .Y(_7860_) );
NOR2X1 NOR2X1_568 ( .gnd(gnd), .vdd(vdd), .A(_7577_), .B(_7859_), .Y(_7861_) );
INVX1 INVX1_1047 ( .gnd(gnd), .vdd(vdd), .A(_7861_), .Y(_7862_) );
NAND3X1 NAND3X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_7753_), .B(_7860_), .C(_7862_), .Y(_7863_) );
INVX1 INVX1_1048 ( .gnd(gnd), .vdd(vdd), .A(_7860_), .Y(_7864_) );
OAI21X1 OAI21X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_7864_), .B(_7861_), .C(_7610_), .Y(_7865_) );
AOI21X1 AOI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_7865_), .B(_7863_), .C(module_1_W_146_), .Y(_7866_) );
INVX1 INVX1_1049 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_146_), .Y(_7867_) );
NOR3X1 NOR3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_7610_), .B(_7861_), .C(_7864_), .Y(_7868_) );
AOI21X1 AOI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_7860_), .B(_7862_), .C(_7753_), .Y(_7869_) );
NOR3X1 NOR3X1_222 ( .gnd(gnd), .vdd(vdd), .A(_7868_), .B(_7867_), .C(_7869_), .Y(_7870_) );
NOR2X1 NOR2X1_569 ( .gnd(gnd), .vdd(vdd), .A(_7866_), .B(_7870_), .Y(_7871_) );
NAND2X1 NAND2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_7643_), .B(_7871_), .Y(_7872_) );
OAI21X1 OAI21X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_7870_), .B(_7866_), .C(_7654_), .Y(_7873_) );
AND2X2 AND2X2_165 ( .gnd(gnd), .vdd(vdd), .A(_7872_), .B(_7873_), .Y(_7874_) );
NAND2X1 NAND2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_7687_), .B(_7874_), .Y(_7875_) );
INVX1 INVX1_1050 ( .gnd(gnd), .vdd(vdd), .A(_7875_), .Y(_7876_) );
NOR2X1 NOR2X1_570 ( .gnd(gnd), .vdd(vdd), .A(_7687_), .B(_7874_), .Y(_7877_) );
OAI21X1 OAI21X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_7876_), .B(_7877_), .C(_7752_), .Y(_7878_) );
NOR2X1 NOR2X1_571 ( .gnd(gnd), .vdd(vdd), .A(_7877_), .B(_7876_), .Y(_7879_) );
NAND2X1 NAND2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_162_), .B(_7879_), .Y(_7880_) );
NAND3X1 NAND3X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_7707_), .B(_7878_), .C(_7880_), .Y(_7881_) );
INVX1 INVX1_1051 ( .gnd(gnd), .vdd(vdd), .A(_7878_), .Y(_7882_) );
AND2X2 AND2X2_166 ( .gnd(gnd), .vdd(vdd), .A(_7879_), .B(module_1_W_162_), .Y(_7883_) );
OAI21X1 OAI21X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_7883_), .B(_7882_), .C(_7708_), .Y(_7884_) );
NAND3X1 NAND3X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_7711_), .B(_7881_), .C(_7884_), .Y(_7885_) );
INVX2 INVX2_249 ( .gnd(gnd), .vdd(vdd), .A(_7885_), .Y(_7886_) );
AOI21X1 AOI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_7881_), .B(_7884_), .C(_7711_), .Y(_7887_) );
OAI21X1 OAI21X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_7886_), .B(_7887_), .C(_7751_), .Y(_7888_) );
NOR2X1 NOR2X1_572 ( .gnd(gnd), .vdd(vdd), .A(_7887_), .B(_7886_), .Y(_7889_) );
NAND2X1 NAND2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_178_), .B(_7889_), .Y(_7890_) );
NAND3X1 NAND3X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_7717_), .B(_7888_), .C(_7890_), .Y(_7891_) );
INVX1 INVX1_1052 ( .gnd(gnd), .vdd(vdd), .A(_7888_), .Y(_7892_) );
INVX1 INVX1_1053 ( .gnd(gnd), .vdd(vdd), .A(_7890_), .Y(_7893_) );
OAI21X1 OAI21X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_7893_), .B(_7892_), .C(_7716_), .Y(_7894_) );
NAND3X1 NAND3X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_7720_), .B(_7891_), .C(_7894_), .Y(_7895_) );
INVX2 INVX2_250 ( .gnd(gnd), .vdd(vdd), .A(_7895_), .Y(_7896_) );
AOI21X1 AOI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_7891_), .B(_7894_), .C(_7720_), .Y(_7897_) );
OAI21X1 OAI21X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_7896_), .B(_7897_), .C(_7750_), .Y(_7898_) );
INVX1 INVX1_1054 ( .gnd(gnd), .vdd(vdd), .A(_7898_), .Y(_7899_) );
NOR3X1 NOR3X1_223 ( .gnd(gnd), .vdd(vdd), .A(_7750_), .B(_7897_), .C(_7896_), .Y(_7900_) );
NOR2X1 NOR2X1_573 ( .gnd(gnd), .vdd(vdd), .A(_7900_), .B(_7899_), .Y(_7901_) );
NAND2X1 NAND2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_7724_), .B(_7901_), .Y(_7902_) );
OAI21X1 OAI21X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_7899_), .B(_7900_), .C(_7725_), .Y(_7903_) );
NAND3X1 NAND3X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_7728_), .B(_7903_), .C(_7902_), .Y(_7904_) );
INVX2 INVX2_251 ( .gnd(gnd), .vdd(vdd), .A(_7904_), .Y(_7905_) );
AOI21X1 AOI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_7903_), .B(_7902_), .C(_7728_), .Y(_7906_) );
NOR2X1 NOR2X1_574 ( .gnd(gnd), .vdd(vdd), .A(_7906_), .B(_7905_), .Y(_7907_) );
NOR2X1 NOR2X1_575 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_210_), .B(_7907_), .Y(_7908_) );
INVX1 INVX1_1055 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_210_), .Y(_7909_) );
NOR3X1 NOR3X1_224 ( .gnd(gnd), .vdd(vdd), .A(_7909_), .B(_7906_), .C(_7905_), .Y(_7910_) );
NOR2X1 NOR2X1_576 ( .gnd(gnd), .vdd(vdd), .A(_7910_), .B(_7908_), .Y(_7911_) );
NAND2X1 NAND2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_7734_), .B(_7911_), .Y(_7912_) );
INVX1 INVX1_1056 ( .gnd(gnd), .vdd(vdd), .A(_7912_), .Y(_7913_) );
OAI21X1 OAI21X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_7908_), .B(_7910_), .C(_7733_), .Y(_7914_) );
INVX2 INVX2_252 ( .gnd(gnd), .vdd(vdd), .A(_7914_), .Y(_7915_) );
NOR2X1 NOR2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_7915_), .B(_7913_), .Y(_7916_) );
NAND2X1 NAND2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_7737_), .B(_7916_), .Y(_7917_) );
OAI21X1 OAI21X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_7913_), .B(_7915_), .C(_7738_), .Y(_7918_) );
AOI21X1 AOI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_7918_), .B(_7917_), .C(module_1_W_226_), .Y(_7919_) );
INVX1 INVX1_1057 ( .gnd(gnd), .vdd(vdd), .A(_7919_), .Y(_7920_) );
NAND3X1 NAND3X1_1801 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_226_), .B(_7918_), .C(_7917_), .Y(_7921_) );
NAND3X1 NAND3X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_7741_), .B(_7921_), .C(_7920_), .Y(_7922_) );
INVX2 INVX2_253 ( .gnd(gnd), .vdd(vdd), .A(_7921_), .Y(_7923_) );
OAI21X1 OAI21X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_7923_), .B(_7919_), .C(_7742_), .Y(_7924_) );
NAND3X1 NAND3X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_7745_), .B(_7924_), .C(_7922_), .Y(_7925_) );
INVX1 INVX1_1058 ( .gnd(gnd), .vdd(vdd), .A(_7925_), .Y(_7926_) );
AOI21X1 AOI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_7924_), .B(_7922_), .C(_7745_), .Y(_7927_) );
OAI21X1 OAI21X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_7926_), .B(_7927_), .C(_7749_), .Y(_7928_) );
NOR2X1 NOR2X1_578 ( .gnd(gnd), .vdd(vdd), .A(_7927_), .B(_7926_), .Y(_7929_) );
NAND2X1 NAND2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_242_), .B(_7929_), .Y(_7930_) );
NAND3X1 NAND3X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_7748_), .B(_7928_), .C(_7930_), .Y(_7931_) );
NAND2X1 NAND2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_224_), .B(_6689_), .Y(_7932_) );
OR2X2 OR2X2_172 ( .gnd(gnd), .vdd(vdd), .A(_6689_), .B(module_1_W_224_), .Y(_7933_) );
NAND2X1 NAND2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_7932_), .B(_7933_), .Y(_7934_) );
INVX4 INVX4_6 ( .gnd(gnd), .vdd(vdd), .A(_7934_), .Y(_7935_) );
INVX2 INVX2_254 ( .gnd(gnd), .vdd(vdd), .A(_7747_), .Y(_7936_) );
NOR2X1 NOR2X1_579 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_241_), .B(_7936_), .Y(_7937_) );
NOR2X1 NOR2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_7748_), .B(_7937_), .Y(_7938_) );
OAI21X1 OAI21X1_1239 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_240_), .B(_7935_), .C(_7938_), .Y(_7939_) );
INVX1 INVX1_1059 ( .gnd(gnd), .vdd(vdd), .A(_7748_), .Y(_7940_) );
INVX1 INVX1_1060 ( .gnd(gnd), .vdd(vdd), .A(_7928_), .Y(_7941_) );
INVX1 INVX1_1061 ( .gnd(gnd), .vdd(vdd), .A(_7930_), .Y(_7942_) );
OAI21X1 OAI21X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_7942_), .B(_7941_), .C(_7940_), .Y(_7943_) );
INVX1 INVX1_1062 ( .gnd(gnd), .vdd(vdd), .A(_7943_), .Y(_7944_) );
OAI21X1 OAI21X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_7944_), .B(_7939_), .C(_7931_), .Y(_7945_) );
INVX1 INVX1_1063 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_243_), .Y(_7946_) );
NAND2X1 NAND2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_7922_), .B(_7925_), .Y(_7947_) );
INVX1 INVX1_1064 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_227_), .Y(_7948_) );
OAI21X1 OAI21X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_7738_), .B(_7915_), .C(_7912_), .Y(_7949_) );
INVX1 INVX1_1065 ( .gnd(gnd), .vdd(vdd), .A(_7910_), .Y(_7950_) );
INVX1 INVX1_1066 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_211_), .Y(_7951_) );
INVX1 INVX1_1067 ( .gnd(gnd), .vdd(vdd), .A(_7902_), .Y(_7952_) );
AOI21X1 AOI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_7728_), .B(_7903_), .C(_7952_), .Y(_7953_) );
INVX1 INVX1_1068 ( .gnd(gnd), .vdd(vdd), .A(_7900_), .Y(_7954_) );
INVX1 INVX1_1069 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_195_), .Y(_7955_) );
AND2X2 AND2X2_167 ( .gnd(gnd), .vdd(vdd), .A(_7895_), .B(_7891_), .Y(_7956_) );
INVX1 INVX1_1070 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_179_), .Y(_7957_) );
INVX1 INVX1_1071 ( .gnd(gnd), .vdd(vdd), .A(_7881_), .Y(_7958_) );
INVX1 INVX1_1072 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_163_), .Y(_7959_) );
INVX1 INVX1_1073 ( .gnd(gnd), .vdd(vdd), .A(_7873_), .Y(_7960_) );
OAI21X1 OAI21X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_7698_), .B(_7960_), .C(_7872_), .Y(_7961_) );
INVX1 INVX1_1074 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_147_), .Y(_7962_) );
OAI21X1 OAI21X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_7610_), .B(_7861_), .C(_7860_), .Y(_7963_) );
INVX1 INVX1_1075 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_131_), .Y(_7964_) );
OAI21X1 OAI21X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_7533_), .B(_7852_), .C(_7848_), .Y(_7965_) );
OAI21X1 OAI21X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_7840_), .B(_7838_), .C(_7832_), .Y(_7966_) );
OAI21X1 OAI21X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_7829_), .B(_7827_), .C(_7821_), .Y(_7967_) );
INVX1 INVX1_1076 ( .gnd(gnd), .vdd(vdd), .A(_7819_), .Y(_7968_) );
AND2X2 AND2X2_168 ( .gnd(gnd), .vdd(vdd), .A(_7813_), .B(_7809_), .Y(_7969_) );
AOI21X1 AOI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_7803_), .B(_7237_), .C(_7796_), .Y(_7970_) );
INVX2 INVX2_255 ( .gnd(gnd), .vdd(vdd), .A(_7970_), .Y(_7971_) );
OAI21X1 OAI21X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_7793_), .B(_7791_), .C(_7782_), .Y(_7972_) );
NOR3X1 NOR3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_7771_), .B(_7138_), .C(_7772_), .Y(_7973_) );
AOI21X1 AOI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_7776_), .B(_7773_), .C(_7973_), .Y(_7974_) );
INVX1 INVX1_1077 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_19_), .Y(_7975_) );
INVX2 INVX2_256 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_3_), .Y(_7976_) );
NOR2X1 NOR2X1_581 ( .gnd(gnd), .vdd(vdd), .A(_7976_), .B(_7764_), .Y(_7977_) );
AND2X2 AND2X2_169 ( .gnd(gnd), .vdd(vdd), .A(_7764_), .B(_7976_), .Y(_7978_) );
OAI21X1 OAI21X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_7978_), .B(_7977_), .C(_7975_), .Y(_7979_) );
NOR2X1 NOR2X1_582 ( .gnd(gnd), .vdd(vdd), .A(_7977_), .B(_7978_), .Y(_7980_) );
NAND2X1 NAND2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_19_), .B(_7980_), .Y(_7981_) );
AOI21X1 AOI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_7979_), .B(_7981_), .C(_7769_), .Y(_7982_) );
INVX1 INVX1_1078 ( .gnd(gnd), .vdd(vdd), .A(_7977_), .Y(_7983_) );
NAND2X1 NAND2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_7976_), .B(_7764_), .Y(_7984_) );
AOI21X1 AOI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_7984_), .B(_7983_), .C(module_1_W_19_), .Y(_7985_) );
NOR3X1 NOR3X1_226 ( .gnd(gnd), .vdd(vdd), .A(_7977_), .B(_7975_), .C(_7978_), .Y(_7986_) );
NOR3X1 NOR3X1_227 ( .gnd(gnd), .vdd(vdd), .A(_7772_), .B(_7986_), .C(_7985_), .Y(_7987_) );
OAI21X1 OAI21X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_7982_), .B(_7987_), .C(_7974_), .Y(_7988_) );
NOR2X1 NOR2X1_583 ( .gnd(gnd), .vdd(vdd), .A(_7987_), .B(_7982_), .Y(_7989_) );
OAI21X1 OAI21X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_7775_), .B(_7973_), .C(_7989_), .Y(_7990_) );
AOI21X1 AOI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_7988_), .B(_7990_), .C(bloque_datos_3_bF_buf3_), .Y(_7991_) );
INVX1 INVX1_1079 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf2_), .Y(_7992_) );
INVX1 INVX1_1080 ( .gnd(gnd), .vdd(vdd), .A(_7988_), .Y(_7993_) );
AOI21X1 AOI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_7769_), .B(_7767_), .C(_7095_), .Y(_7994_) );
OAI21X1 OAI21X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_7994_), .B(_7149_), .C(_7770_), .Y(_7995_) );
AND2X2 AND2X2_170 ( .gnd(gnd), .vdd(vdd), .A(_7989_), .B(_7995_), .Y(_7996_) );
NOR3X1 NOR3X1_228 ( .gnd(gnd), .vdd(vdd), .A(_7993_), .B(_7992_), .C(_7996_), .Y(_7997_) );
OAI21X1 OAI21X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_7997_), .B(_7991_), .C(_7784_), .Y(_7998_) );
OAI21X1 OAI21X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_7996_), .B(_7993_), .C(_7992_), .Y(_7999_) );
NAND3X1 NAND3X1_1805 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf1_), .B(_7988_), .C(_7990_), .Y(_8000_) );
NAND3X1 NAND3X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_7781_), .B(_8000_), .C(_7999_), .Y(_8001_) );
AOI21X1 AOI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_8001_), .B(_7998_), .C(_7972_), .Y(_8002_) );
INVX2 INVX2_257 ( .gnd(gnd), .vdd(vdd), .A(_8002_), .Y(_8003_) );
NAND3X1 NAND3X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_7972_), .B(_8001_), .C(_7998_), .Y(_8004_) );
AOI21X1 AOI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_8004_), .B(_8003_), .C(bloque_datos_19_bF_buf3_), .Y(_8005_) );
INVX1 INVX1_1081 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf2_), .Y(_8006_) );
INVX2 INVX2_258 ( .gnd(gnd), .vdd(vdd), .A(_8004_), .Y(_8007_) );
NOR3X1 NOR3X1_229 ( .gnd(gnd), .vdd(vdd), .A(_8006_), .B(_8002_), .C(_8007_), .Y(_8008_) );
OAI21X1 OAI21X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_8008_), .B(_8005_), .C(_7795_), .Y(_8009_) );
OAI21X1 OAI21X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_8007_), .B(_8002_), .C(_8006_), .Y(_8010_) );
NAND3X1 NAND3X1_1808 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf1_), .B(_8004_), .C(_8003_), .Y(_8011_) );
NAND3X1 NAND3X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_7799_), .B(_8010_), .C(_8011_), .Y(_8012_) );
AOI21X1 AOI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_8012_), .B(_8009_), .C(_7971_), .Y(_8013_) );
NAND2X1 NAND2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_8012_), .B(_8009_), .Y(_8014_) );
NOR2X1 NOR2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_7970_), .B(_8014_), .Y(_8015_) );
OAI21X1 OAI21X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_8015_), .B(_8013_), .C(bloque_datos_35_bF_buf3_), .Y(_8016_) );
INVX1 INVX1_1082 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf2_), .Y(_8017_) );
INVX1 INVX1_1083 ( .gnd(gnd), .vdd(vdd), .A(_8009_), .Y(_8018_) );
INVX1 INVX1_1084 ( .gnd(gnd), .vdd(vdd), .A(_8012_), .Y(_8019_) );
OAI21X1 OAI21X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_8018_), .B(_8019_), .C(_7970_), .Y(_8020_) );
NAND3X1 NAND3X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_8012_), .B(_8009_), .C(_7971_), .Y(_8021_) );
NAND3X1 NAND3X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_8017_), .B(_8021_), .C(_8020_), .Y(_8022_) );
NAND3X1 NAND3X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_7811_), .B(_8022_), .C(_8016_), .Y(_8023_) );
OAI21X1 OAI21X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_8015_), .B(_8013_), .C(_8017_), .Y(_8024_) );
NAND3X1 NAND3X1_1813 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf1_), .B(_8021_), .C(_8020_), .Y(_8025_) );
NAND3X1 NAND3X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_7808_), .B(_8025_), .C(_8024_), .Y(_8026_) );
NAND2X1 NAND2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_8023_), .B(_8026_), .Y(_8027_) );
NAND2X1 NAND2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_8027_), .B(_7969_), .Y(_8028_) );
OR2X2 OR2X2_173 ( .gnd(gnd), .vdd(vdd), .A(_7969_), .B(_8027_), .Y(_8029_) );
NAND2X1 NAND2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_8028_), .B(_8029_), .Y(_8030_) );
XNOR2X1 XNOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_8030_), .B(bloque_datos_51_bF_buf3_), .Y(_8031_) );
OR2X2 OR2X2_174 ( .gnd(gnd), .vdd(vdd), .A(_8031_), .B(_7968_), .Y(_8032_) );
NOR2X1 NOR2X1_585 ( .gnd(gnd), .vdd(vdd), .A(_7814_), .B(_7818_), .Y(_8033_) );
INVX2 INVX2_259 ( .gnd(gnd), .vdd(vdd), .A(_8033_), .Y(_8034_) );
OAI21X1 OAI21X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_7817_), .B(_8034_), .C(_8031_), .Y(_8035_) );
AOI21X1 AOI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_8035_), .B(_8032_), .C(_7967_), .Y(_8036_) );
INVX2 INVX2_260 ( .gnd(gnd), .vdd(vdd), .A(_7967_), .Y(_8037_) );
NOR2X1 NOR2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_7968_), .B(_8031_), .Y(_8038_) );
NAND2X1 NAND2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf2_), .B(_8030_), .Y(_8039_) );
OR2X2 OR2X2_175 ( .gnd(gnd), .vdd(vdd), .A(_8030_), .B(bloque_datos_51_bF_buf1_), .Y(_8040_) );
AOI21X1 AOI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_8039_), .B(_8040_), .C(_7819_), .Y(_8041_) );
NOR3X1 NOR3X1_230 ( .gnd(gnd), .vdd(vdd), .A(_8037_), .B(_8041_), .C(_8038_), .Y(_8042_) );
OAI21X1 OAI21X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_8036_), .B(_8042_), .C(bloque_datos_67_bF_buf2_), .Y(_8043_) );
INVX1 INVX1_1085 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf1_), .Y(_8044_) );
NOR2X1 NOR2X1_587 ( .gnd(gnd), .vdd(vdd), .A(_8042_), .B(_8036_), .Y(_8045_) );
NAND2X1 NAND2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_8044_), .B(_8045_), .Y(_8046_) );
NAND3X1 NAND3X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_7835_), .B(_8043_), .C(_8046_), .Y(_8047_) );
OAI21X1 OAI21X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_8036_), .B(_8042_), .C(_8044_), .Y(_8048_) );
NAND2X1 NAND2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf0_), .B(_8045_), .Y(_8049_) );
NAND3X1 NAND3X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_7831_), .B(_8048_), .C(_8049_), .Y(_8050_) );
AOI21X1 AOI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_8050_), .B(_8047_), .C(_7966_), .Y(_8051_) );
NAND3X1 NAND3X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_7966_), .B(_8050_), .C(_8047_), .Y(_8052_) );
INVX2 INVX2_261 ( .gnd(gnd), .vdd(vdd), .A(_8052_), .Y(_8053_) );
OAI21X1 OAI21X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_8053_), .B(_8051_), .C(bloque_datos_83_bF_buf3_), .Y(_8054_) );
INVX1 INVX1_1086 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf2_), .Y(_8055_) );
INVX2 INVX2_262 ( .gnd(gnd), .vdd(vdd), .A(_8051_), .Y(_8056_) );
NAND3X1 NAND3X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_8055_), .B(_8052_), .C(_8056_), .Y(_8057_) );
NAND3X1 NAND3X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_7846_), .B(_8057_), .C(_8054_), .Y(_8058_) );
INVX1 INVX1_1087 ( .gnd(gnd), .vdd(vdd), .A(_7846_), .Y(_8059_) );
OAI21X1 OAI21X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_8053_), .B(_8051_), .C(_8055_), .Y(_8060_) );
NAND3X1 NAND3X1_1820 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf1_), .B(_8052_), .C(_8056_), .Y(_8061_) );
NAND3X1 NAND3X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_8059_), .B(_8061_), .C(_8060_), .Y(_8062_) );
AOI21X1 AOI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_8058_), .B(_8062_), .C(_7965_), .Y(_8063_) );
NAND3X1 NAND3X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_7965_), .B(_8058_), .C(_8062_), .Y(_8064_) );
INVX2 INVX2_263 ( .gnd(gnd), .vdd(vdd), .A(_8064_), .Y(_8065_) );
OAI21X1 OAI21X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_8065_), .B(_8063_), .C(_7964_), .Y(_8066_) );
INVX1 INVX1_1088 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .Y(_8067_) );
NAND3X1 NAND3X1_1823 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_131_), .B(_8064_), .C(_8067_), .Y(_8068_) );
NAND2X1 NAND2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_8068_), .B(_8066_), .Y(_8069_) );
NAND2X1 NAND2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_7858_), .B(_8069_), .Y(_8070_) );
INVX1 INVX1_1089 ( .gnd(gnd), .vdd(vdd), .A(_7858_), .Y(_8071_) );
NAND3X1 NAND3X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_8071_), .B(_8068_), .C(_8066_), .Y(_8072_) );
NAND3X1 NAND3X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_8072_), .B(_8070_), .C(_7963_), .Y(_8073_) );
INVX1 INVX1_1090 ( .gnd(gnd), .vdd(vdd), .A(_8073_), .Y(_8074_) );
AND2X2 AND2X2_171 ( .gnd(gnd), .vdd(vdd), .A(_8070_), .B(_8072_), .Y(_8075_) );
NOR2X1 NOR2X1_588 ( .gnd(gnd), .vdd(vdd), .A(_7963_), .B(_8075_), .Y(_8076_) );
OAI21X1 OAI21X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_8076_), .B(_8074_), .C(_7962_), .Y(_8077_) );
NOR3X1 NOR3X1_231 ( .gnd(gnd), .vdd(vdd), .A(_7962_), .B(_8074_), .C(_8076_), .Y(_8078_) );
INVX2 INVX2_264 ( .gnd(gnd), .vdd(vdd), .A(_8078_), .Y(_8079_) );
NAND3X1 NAND3X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_7870_), .B(_8077_), .C(_8079_), .Y(_8080_) );
INVX1 INVX1_1091 ( .gnd(gnd), .vdd(vdd), .A(_7870_), .Y(_8081_) );
INVX1 INVX1_1092 ( .gnd(gnd), .vdd(vdd), .A(_8077_), .Y(_8082_) );
OAI21X1 OAI21X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_8082_), .B(_8078_), .C(_8081_), .Y(_8083_) );
NAND3X1 NAND3X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_8083_), .B(_7961_), .C(_8080_), .Y(_8084_) );
INVX1 INVX1_1093 ( .gnd(gnd), .vdd(vdd), .A(_8084_), .Y(_8085_) );
AOI21X1 AOI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_8083_), .B(_8080_), .C(_7961_), .Y(_8086_) );
OAI21X1 OAI21X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_8085_), .B(_8086_), .C(_7959_), .Y(_8087_) );
NOR2X1 NOR2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_8086_), .B(_8085_), .Y(_8088_) );
NAND2X1 NAND2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_163_), .B(_8088_), .Y(_8089_) );
NAND2X1 NAND2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_8087_), .B(_8089_), .Y(_8090_) );
NOR2X1 NOR2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_7880_), .B(_8090_), .Y(_8091_) );
INVX2 INVX2_265 ( .gnd(gnd), .vdd(vdd), .A(_7879_), .Y(_8092_) );
OAI21X1 OAI21X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_7752_), .B(_8092_), .C(_8090_), .Y(_8093_) );
INVX2 INVX2_266 ( .gnd(gnd), .vdd(vdd), .A(_8093_), .Y(_8094_) );
NOR2X1 NOR2X1_591 ( .gnd(gnd), .vdd(vdd), .A(_8091_), .B(_8094_), .Y(_8095_) );
OAI21X1 OAI21X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_7886_), .B(_7958_), .C(_8095_), .Y(_8096_) );
AOI21X1 AOI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_7711_), .B(_7884_), .C(_7958_), .Y(_8097_) );
OAI21X1 OAI21X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_8094_), .B(_8091_), .C(_8097_), .Y(_8098_) );
NAND2X1 NAND2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_8098_), .B(_8096_), .Y(_8099_) );
NAND2X1 NAND2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_7957_), .B(_8099_), .Y(_8100_) );
NOR2X1 NOR2X1_592 ( .gnd(gnd), .vdd(vdd), .A(_7957_), .B(_8099_), .Y(_8101_) );
INVX2 INVX2_267 ( .gnd(gnd), .vdd(vdd), .A(_8101_), .Y(_8102_) );
NAND3X1 NAND3X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_7893_), .B(_8100_), .C(_8102_), .Y(_8103_) );
INVX1 INVX1_1094 ( .gnd(gnd), .vdd(vdd), .A(_8100_), .Y(_8104_) );
OAI21X1 OAI21X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_8104_), .B(_8101_), .C(_7890_), .Y(_8105_) );
NAND2X1 NAND2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_8105_), .B(_8103_), .Y(_8106_) );
NOR2X1 NOR2X1_593 ( .gnd(gnd), .vdd(vdd), .A(_7956_), .B(_8106_), .Y(_8107_) );
INVX1 INVX1_1095 ( .gnd(gnd), .vdd(vdd), .A(_8103_), .Y(_8108_) );
INVX1 INVX1_1096 ( .gnd(gnd), .vdd(vdd), .A(_8105_), .Y(_8109_) );
OAI21X1 OAI21X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_8108_), .B(_8109_), .C(_7956_), .Y(_8110_) );
INVX1 INVX1_1097 ( .gnd(gnd), .vdd(vdd), .A(_8110_), .Y(_8111_) );
OAI21X1 OAI21X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_8111_), .B(_8107_), .C(_7955_), .Y(_8112_) );
NOR2X1 NOR2X1_594 ( .gnd(gnd), .vdd(vdd), .A(_8107_), .B(_8111_), .Y(_8113_) );
NAND2X1 NAND2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_195_), .B(_8113_), .Y(_8114_) );
NAND2X1 NAND2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_8112_), .B(_8114_), .Y(_8115_) );
OR2X2 OR2X2_176 ( .gnd(gnd), .vdd(vdd), .A(_8115_), .B(_7954_), .Y(_8116_) );
AOI21X1 AOI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_8112_), .B(_8114_), .C(_7900_), .Y(_8117_) );
INVX1 INVX1_1098 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .Y(_8118_) );
NAND2X1 NAND2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_8118_), .B(_8116_), .Y(_8119_) );
NOR2X1 NOR2X1_595 ( .gnd(gnd), .vdd(vdd), .A(_7953_), .B(_8119_), .Y(_8120_) );
NOR2X1 NOR2X1_596 ( .gnd(gnd), .vdd(vdd), .A(_7954_), .B(_8115_), .Y(_8121_) );
OAI21X1 OAI21X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_8121_), .B(_8117_), .C(_7953_), .Y(_8122_) );
INVX2 INVX2_268 ( .gnd(gnd), .vdd(vdd), .A(_8122_), .Y(_8123_) );
OAI21X1 OAI21X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_8120_), .B(_8123_), .C(_7951_), .Y(_8124_) );
INVX1 INVX1_1099 ( .gnd(gnd), .vdd(vdd), .A(_8124_), .Y(_8125_) );
NOR2X1 NOR2X1_597 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .B(_8121_), .Y(_8126_) );
OAI21X1 OAI21X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_7952_), .B(_7905_), .C(_8126_), .Y(_8127_) );
NAND2X1 NAND2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_8122_), .B(_8127_), .Y(_8128_) );
NOR2X1 NOR2X1_598 ( .gnd(gnd), .vdd(vdd), .A(_7951_), .B(_8128_), .Y(_8129_) );
NOR3X1 NOR3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_7950_), .B(_8129_), .C(_8125_), .Y(_8130_) );
NOR2X1 NOR2X1_599 ( .gnd(gnd), .vdd(vdd), .A(_8123_), .B(_8120_), .Y(_8131_) );
NAND2X1 NAND2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_211_), .B(_8131_), .Y(_8132_) );
AOI21X1 AOI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_8124_), .B(_8132_), .C(_7910_), .Y(_8133_) );
NOR2X1 NOR2X1_600 ( .gnd(gnd), .vdd(vdd), .A(_8133_), .B(_8130_), .Y(_8134_) );
AND2X2 AND2X2_172 ( .gnd(gnd), .vdd(vdd), .A(_8134_), .B(_7949_), .Y(_8135_) );
INVX1 INVX1_1100 ( .gnd(gnd), .vdd(vdd), .A(_7949_), .Y(_8136_) );
OAI21X1 OAI21X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_8130_), .B(_8133_), .C(_8136_), .Y(_8137_) );
INVX2 INVX2_269 ( .gnd(gnd), .vdd(vdd), .A(_8137_), .Y(_8138_) );
OAI21X1 OAI21X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_8135_), .B(_8138_), .C(_7948_), .Y(_8139_) );
NOR2X1 NOR2X1_601 ( .gnd(gnd), .vdd(vdd), .A(_8138_), .B(_8135_), .Y(_8140_) );
NAND2X1 NAND2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_227_), .B(_8140_), .Y(_8141_) );
NAND3X1 NAND3X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_7923_), .B(_8139_), .C(_8141_), .Y(_8142_) );
NAND2X1 NAND2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_8139_), .B(_8141_), .Y(_8143_) );
NAND2X1 NAND2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_7921_), .B(_8143_), .Y(_8144_) );
NAND3X1 NAND3X1_1830 ( .gnd(gnd), .vdd(vdd), .A(_7947_), .B(_8142_), .C(_8144_), .Y(_8145_) );
INVX2 INVX2_270 ( .gnd(gnd), .vdd(vdd), .A(_8145_), .Y(_8146_) );
AND2X2 AND2X2_173 ( .gnd(gnd), .vdd(vdd), .A(_7925_), .B(_7922_), .Y(_8147_) );
INVX1 INVX1_1101 ( .gnd(gnd), .vdd(vdd), .A(_8142_), .Y(_8148_) );
AOI21X1 AOI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_8139_), .B(_8141_), .C(_7923_), .Y(_8149_) );
OAI21X1 OAI21X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_8148_), .B(_8149_), .C(_8147_), .Y(_8150_) );
INVX2 INVX2_271 ( .gnd(gnd), .vdd(vdd), .A(_8150_), .Y(_8151_) );
OAI21X1 OAI21X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_8151_), .B(_8146_), .C(_7946_), .Y(_8152_) );
NOR2X1 NOR2X1_602 ( .gnd(gnd), .vdd(vdd), .A(_8146_), .B(_8151_), .Y(_8153_) );
NAND2X1 NAND2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_243_), .B(_8153_), .Y(_8154_) );
NAND2X1 NAND2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_8152_), .B(_8154_), .Y(_8155_) );
OR2X2 OR2X2_177 ( .gnd(gnd), .vdd(vdd), .A(_8155_), .B(_7930_), .Y(_8156_) );
INVX2 INVX2_272 ( .gnd(gnd), .vdd(vdd), .A(_7929_), .Y(_8157_) );
OAI21X1 OAI21X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_8157_), .B(_7749_), .C(_8155_), .Y(_8158_) );
AOI21X1 AOI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_8158_), .B(_8156_), .C(_7945_), .Y(_8159_) );
INVX1 INVX1_1102 ( .gnd(gnd), .vdd(vdd), .A(_7945_), .Y(_8160_) );
NAND2X1 NAND2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_8158_), .B(_8156_), .Y(_8161_) );
NOR2X1 NOR2X1_603 ( .gnd(gnd), .vdd(vdd), .A(_8160_), .B(_8161_), .Y(_8162_) );
NOR2X1 NOR2X1_604 ( .gnd(gnd), .vdd(vdd), .A(_8159_), .B(_8162_), .Y(_8163_) );
INVX2 INVX2_273 ( .gnd(gnd), .vdd(vdd), .A(_8163_), .Y(module_1_H_15_) );
NOR2X1 NOR2X1_605 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_240_), .B(_7935_), .Y(_8164_) );
OAI21X1 OAI21X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_7937_), .B(_7748_), .C(_8164_), .Y(_8165_) );
NAND2X1 NAND2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_8165_), .B(_7939_), .Y(_8166_) );
INVX2 INVX2_274 ( .gnd(gnd), .vdd(vdd), .A(_8166_), .Y(module_1_H_13_) );
NAND2X1 NAND2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_240_), .B(_7935_), .Y(_8167_) );
INVX1 INVX1_1103 ( .gnd(gnd), .vdd(vdd), .A(_8167_), .Y(_8168_) );
NOR2X1 NOR2X1_606 ( .gnd(gnd), .vdd(vdd), .A(_8164_), .B(_8168_), .Y(module_1_H_0_) );
INVX1 INVX1_1104 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_0_), .Y(module_1_H_12_) );
INVX1 INVX1_1105 ( .gnd(gnd), .vdd(vdd), .A(_7939_), .Y(_8169_) );
OAI21X1 OAI21X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_8164_), .B(_8168_), .C(module_1_H_13_), .Y(_8170_) );
INVX2 INVX2_275 ( .gnd(gnd), .vdd(vdd), .A(_8170_), .Y(_8171_) );
AOI21X1 AOI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_8169_), .B(_8167_), .C(_8171_), .Y(module_1_H_1_) );
NAND3X1 NAND3X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_7931_), .B(_8169_), .C(_7943_), .Y(_8172_) );
INVX1 INVX1_1106 ( .gnd(gnd), .vdd(vdd), .A(_7931_), .Y(_8173_) );
OAI21X1 OAI21X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_7944_), .B(_8173_), .C(_7939_), .Y(_8174_) );
AND2X2 AND2X2_174 ( .gnd(gnd), .vdd(vdd), .A(_8174_), .B(_8172_), .Y(module_1_H_14_) );
NAND2X1 NAND2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_8171_), .B(module_1_H_14_), .Y(_8175_) );
INVX1 INVX1_1107 ( .gnd(gnd), .vdd(vdd), .A(_8175_), .Y(_8176_) );
NOR2X1 NOR2X1_607 ( .gnd(gnd), .vdd(vdd), .A(_8171_), .B(module_1_H_14_), .Y(_8177_) );
NOR2X1 NOR2X1_608 ( .gnd(gnd), .vdd(vdd), .A(_8177_), .B(_8176_), .Y(module_1_H_2_) );
NOR3X1 NOR3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_8175_), .B(_8159_), .C(_8162_), .Y(_8178_) );
NOR2X1 NOR2X1_609 ( .gnd(gnd), .vdd(vdd), .A(_8176_), .B(_8163_), .Y(_8179_) );
NOR2X1 NOR2X1_610 ( .gnd(gnd), .vdd(vdd), .A(_8178_), .B(_8179_), .Y(module_1_H_3_) );
AOI21X1 AOI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_8152_), .B(_8154_), .C(_7942_), .Y(_8180_) );
OAI21X1 OAI21X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_8160_), .B(_8180_), .C(_8156_), .Y(_8181_) );
INVX1 INVX1_1108 ( .gnd(gnd), .vdd(vdd), .A(_8154_), .Y(_8182_) );
AOI21X1 AOI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_7947_), .B(_8144_), .C(_8148_), .Y(_8183_) );
OAI21X1 OAI21X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_8125_), .B(_8129_), .C(_7950_), .Y(_8184_) );
AOI21X1 AOI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_7949_), .B(_8184_), .C(_8130_), .Y(_8185_) );
INVX1 INVX1_1109 ( .gnd(gnd), .vdd(vdd), .A(_7953_), .Y(_8186_) );
AOI21X1 AOI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_8186_), .B(_8118_), .C(_8121_), .Y(_8187_) );
NAND2X1 NAND2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_7891_), .B(_7895_), .Y(_8188_) );
AOI21X1 AOI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_8188_), .B(_8105_), .C(_8108_), .Y(_8189_) );
INVX1 INVX1_1110 ( .gnd(gnd), .vdd(vdd), .A(_8091_), .Y(_8190_) );
OAI21X1 OAI21X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_8094_), .B(_8097_), .C(_8190_), .Y(_8191_) );
INVX1 INVX1_1111 ( .gnd(gnd), .vdd(vdd), .A(_8191_), .Y(_8192_) );
AND2X2 AND2X2_175 ( .gnd(gnd), .vdd(vdd), .A(_8084_), .B(_8080_), .Y(_8193_) );
NAND2X1 NAND2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_8070_), .B(_8073_), .Y(_8194_) );
AND2X2 AND2X2_176 ( .gnd(gnd), .vdd(vdd), .A(_8064_), .B(_8058_), .Y(_8195_) );
INVX2 INVX2_276 ( .gnd(gnd), .vdd(vdd), .A(_8060_), .Y(_8196_) );
AOI21X1 AOI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_8048_), .B(_8049_), .C(_7831_), .Y(_8197_) );
AOI21X1 AOI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_7966_), .B(_8050_), .C(_8197_), .Y(_8198_) );
INVX2 INVX2_277 ( .gnd(gnd), .vdd(vdd), .A(_8048_), .Y(_8199_) );
AOI21X1 AOI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_7967_), .B(_8035_), .C(_8038_), .Y(_8200_) );
INVX1 INVX1_1112 ( .gnd(gnd), .vdd(vdd), .A(_8030_), .Y(_8201_) );
NOR2X1 NOR2X1_611 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf0_), .B(_8201_), .Y(_8202_) );
NAND2X1 NAND2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_7809_), .B(_7813_), .Y(_8203_) );
INVX1 INVX1_1113 ( .gnd(gnd), .vdd(vdd), .A(_8023_), .Y(_8204_) );
AOI21X1 AOI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_8026_), .B(_8203_), .C(_8204_), .Y(_8205_) );
INVX2 INVX2_278 ( .gnd(gnd), .vdd(vdd), .A(_8024_), .Y(_8206_) );
AOI21X1 AOI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_8012_), .B(_7971_), .C(_8018_), .Y(_8207_) );
AOI21X1 AOI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_8000_), .B(_7999_), .C(_7781_), .Y(_8208_) );
AOI21X1 AOI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_8001_), .B(_7972_), .C(_8208_), .Y(_8209_) );
OAI21X1 OAI21X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_7985_), .B(_7986_), .C(_7772_), .Y(_8210_) );
OAI21X1 OAI21X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_7974_), .B(_7987_), .C(_8210_), .Y(_8211_) );
INVX1 INVX1_1114 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_4_), .Y(_8212_) );
OAI21X1 OAI21X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_7764_), .B(_7976_), .C(_8212_), .Y(_8213_) );
NAND2X1 NAND2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_4_), .B(_7977_), .Y(_8214_) );
AOI21X1 AOI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_8213_), .B(_8214_), .C(_7007_), .Y(_8215_) );
INVX1 INVX1_1115 ( .gnd(gnd), .vdd(vdd), .A(_8213_), .Y(_8216_) );
NOR3X1 NOR3X1_234 ( .gnd(gnd), .vdd(vdd), .A(_7976_), .B(_8212_), .C(_7764_), .Y(_8217_) );
NOR3X1 NOR3X1_235 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_0_), .B(_8217_), .C(_8216_), .Y(_8218_) );
OAI21X1 OAI21X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_8218_), .B(_8215_), .C(module_1_W_20_), .Y(_8219_) );
INVX1 INVX1_1116 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_20_), .Y(_8220_) );
OAI21X1 OAI21X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_8216_), .B(_8217_), .C(module_1_W_0_), .Y(_8221_) );
NAND3X1 NAND3X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_7007_), .B(_8213_), .C(_8214_), .Y(_8222_) );
NAND3X1 NAND3X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_8220_), .B(_8222_), .C(_8221_), .Y(_8223_) );
NAND3X1 NAND3X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_7979_), .B(_8223_), .C(_8219_), .Y(_8224_) );
OAI21X1 OAI21X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_8218_), .B(_8215_), .C(_8220_), .Y(_8225_) );
NAND3X1 NAND3X1_1835 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_20_), .B(_8222_), .C(_8221_), .Y(_8226_) );
NAND3X1 NAND3X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_7985_), .B(_8226_), .C(_8225_), .Y(_8227_) );
NAND3X1 NAND3X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_8224_), .B(_8227_), .C(_8211_), .Y(_8228_) );
NAND3X1 NAND3X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_7769_), .B(_7979_), .C(_7981_), .Y(_8229_) );
AOI21X1 AOI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_8229_), .B(_7995_), .C(_7982_), .Y(_8230_) );
NAND3X1 NAND3X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_7985_), .B(_8223_), .C(_8219_), .Y(_8231_) );
NAND3X1 NAND3X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_7979_), .B(_8226_), .C(_8225_), .Y(_8232_) );
NAND3X1 NAND3X1_1841 ( .gnd(gnd), .vdd(vdd), .A(_8230_), .B(_8231_), .C(_8232_), .Y(_8233_) );
XNOR2X1 XNOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_6309_), .B(module_1_W_8_), .Y(_8234_) );
INVX1 INVX1_1117 ( .gnd(gnd), .vdd(vdd), .A(_8234_), .Y(_8235_) );
NAND3X1 NAND3X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_8235_), .B(_8233_), .C(_8228_), .Y(_8236_) );
AOI21X1 AOI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_8231_), .B(_8232_), .C(_8230_), .Y(_8237_) );
AOI21X1 AOI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_8224_), .B(_8227_), .C(_8211_), .Y(_8238_) );
OAI21X1 OAI21X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_8237_), .B(_8238_), .C(_8234_), .Y(_8239_) );
AOI21X1 AOI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_8236_), .B(_8239_), .C(bloque_datos_4_bF_buf3_), .Y(_8240_) );
INVX1 INVX1_1118 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf2_), .Y(_8241_) );
NAND3X1 NAND3X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_8234_), .B(_8233_), .C(_8228_), .Y(_8242_) );
OAI21X1 OAI21X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_8237_), .B(_8238_), .C(_8235_), .Y(_8243_) );
AOI21X1 AOI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_8242_), .B(_8243_), .C(_8241_), .Y(_8244_) );
OAI21X1 OAI21X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_8240_), .B(_8244_), .C(_7991_), .Y(_8245_) );
NAND3X1 NAND3X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_8241_), .B(_8242_), .C(_8243_), .Y(_8246_) );
NAND3X1 NAND3X1_1845 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf1_), .B(_8236_), .C(_8239_), .Y(_8247_) );
NAND3X1 NAND3X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_7999_), .B(_8246_), .C(_8247_), .Y(_8248_) );
NAND3X1 NAND3X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_8209_), .B(_8248_), .C(_8245_), .Y(_8249_) );
AOI21X1 AOI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_7785_), .B(_7760_), .C(_7792_), .Y(_8250_) );
NOR3X1 NOR3X1_236 ( .gnd(gnd), .vdd(vdd), .A(_7784_), .B(_7991_), .C(_7997_), .Y(_8251_) );
OAI21X1 OAI21X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_8251_), .B(_8250_), .C(_7998_), .Y(_8252_) );
OAI21X1 OAI21X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_8240_), .B(_8244_), .C(_7999_), .Y(_8253_) );
NAND3X1 NAND3X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_7991_), .B(_8246_), .C(_8247_), .Y(_8254_) );
NAND3X1 NAND3X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_8254_), .B(_8253_), .C(_8252_), .Y(_8255_) );
NOR2X1 NOR2X1_612 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_24_), .B(module_1_W_8_), .Y(_8256_) );
INVX1 INVX1_1119 ( .gnd(gnd), .vdd(vdd), .A(_8256_), .Y(_8257_) );
NAND2X1 NAND2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_24_), .B(module_1_W_8_), .Y(_8258_) );
NAND2X1 NAND2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_8258_), .B(_8257_), .Y(_8259_) );
XNOR2X1 XNOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_6331_), .B(_8259_), .Y(_8260_) );
NAND3X1 NAND3X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_8260_), .B(_8249_), .C(_8255_), .Y(_8261_) );
AOI21X1 AOI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_8254_), .B(_8253_), .C(_8252_), .Y(_8262_) );
AOI21X1 AOI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_8248_), .B(_8245_), .C(_8209_), .Y(_8263_) );
INVX1 INVX1_1120 ( .gnd(gnd), .vdd(vdd), .A(_8260_), .Y(_8264_) );
OAI21X1 OAI21X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_8262_), .B(_8263_), .C(_8264_), .Y(_8265_) );
AOI21X1 AOI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_8261_), .B(_8265_), .C(bloque_datos_20_bF_buf3_), .Y(_8266_) );
INVX1 INVX1_1121 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf2_), .Y(_8267_) );
OAI21X1 OAI21X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_8262_), .B(_8263_), .C(_8260_), .Y(_8268_) );
NAND3X1 NAND3X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_8264_), .B(_8249_), .C(_8255_), .Y(_8269_) );
AOI21X1 AOI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_8269_), .B(_8268_), .C(_8267_), .Y(_8270_) );
OAI21X1 OAI21X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_8266_), .B(_8270_), .C(_8005_), .Y(_8271_) );
NAND3X1 NAND3X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_8267_), .B(_8269_), .C(_8268_), .Y(_8272_) );
NAND3X1 NAND3X1_1853 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf1_), .B(_8261_), .C(_8265_), .Y(_8273_) );
NAND3X1 NAND3X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_8010_), .B(_8272_), .C(_8273_), .Y(_8274_) );
NAND3X1 NAND3X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_8274_), .B(_8271_), .C(_8207_), .Y(_8275_) );
OAI21X1 OAI21X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_8019_), .B(_7970_), .C(_8009_), .Y(_8276_) );
OAI21X1 OAI21X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_8266_), .B(_8270_), .C(_8010_), .Y(_8277_) );
NAND3X1 NAND3X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_8005_), .B(_8272_), .C(_8273_), .Y(_8278_) );
NAND3X1 NAND3X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_8278_), .B(_8276_), .C(_8277_), .Y(_8279_) );
INVX1 INVX1_1122 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .Y(_8280_) );
OR2X2 OR2X2_178 ( .gnd(gnd), .vdd(vdd), .A(_8259_), .B(_8280_), .Y(_8281_) );
NAND2X1 NAND2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_8280_), .B(_8259_), .Y(_8282_) );
NAND2X1 NAND2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_8282_), .B(_8281_), .Y(_8283_) );
INVX2 INVX2_279 ( .gnd(gnd), .vdd(vdd), .A(_8283_), .Y(_8284_) );
XNOR2X1 XNOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_6362_), .B(_8284_), .Y(_8285_) );
NAND3X1 NAND3X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_8285_), .B(_8279_), .C(_8275_), .Y(_8286_) );
AOI21X1 AOI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_8278_), .B(_8277_), .C(_8276_), .Y(_4477_) );
AOI21X1 AOI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_8274_), .B(_8271_), .C(_8207_), .Y(_4478_) );
INVX1 INVX1_1123 ( .gnd(gnd), .vdd(vdd), .A(_8285_), .Y(_4479_) );
OAI21X1 OAI21X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_4477_), .B(_4478_), .C(_4479_), .Y(_4480_) );
AOI21X1 AOI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_8286_), .B(_4480_), .C(bloque_datos_36_bF_buf2_), .Y(_4481_) );
INVX1 INVX1_1124 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf1_), .Y(_4482_) );
NAND3X1 NAND3X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .B(_8279_), .C(_8275_), .Y(_4483_) );
OAI21X1 OAI21X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_4477_), .B(_4478_), .C(_8285_), .Y(_4484_) );
AOI21X1 AOI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_4483_), .B(_4484_), .C(_4482_), .Y(_4485_) );
OAI21X1 OAI21X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_4481_), .B(_4485_), .C(_8206_), .Y(_4486_) );
NAND3X1 NAND3X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4483_), .C(_4484_), .Y(_4487_) );
NAND3X1 NAND3X1_1861 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf0_), .B(_8286_), .C(_4480_), .Y(_4488_) );
NAND3X1 NAND3X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_8024_), .B(_4487_), .C(_4488_), .Y(_4489_) );
NAND3X1 NAND3X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_8205_), .B(_4489_), .C(_4486_), .Y(_4490_) );
OAI21X1 OAI21X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_7969_), .B(_8027_), .C(_8023_), .Y(_4491_) );
OAI21X1 OAI21X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_4481_), .B(_4485_), .C(_8024_), .Y(_4492_) );
NAND3X1 NAND3X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_8206_), .B(_4487_), .C(_4488_), .Y(_4493_) );
NAND3X1 NAND3X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_4491_), .B(_4493_), .C(_4492_), .Y(_4494_) );
NAND2X1 NAND2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf2_), .B(_8283_), .Y(_4495_) );
OR2X2 OR2X2_179 ( .gnd(gnd), .vdd(vdd), .A(_8283_), .B(bloque_datos_24_bF_buf1_), .Y(_4496_) );
NAND2X1 NAND2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_4495_), .B(_4496_), .Y(_4497_) );
INVX2 INVX2_280 ( .gnd(gnd), .vdd(vdd), .A(_4497_), .Y(_4498_) );
XNOR2X1 XNOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_6392_), .B(_4498_), .Y(_4499_) );
NAND3X1 NAND3X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_4499_), .B(_4490_), .C(_4494_), .Y(_4500_) );
AOI21X1 AOI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_4493_), .B(_4492_), .C(_4491_), .Y(_4501_) );
AOI21X1 AOI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_4489_), .B(_4486_), .C(_8205_), .Y(_4502_) );
INVX1 INVX1_1125 ( .gnd(gnd), .vdd(vdd), .A(_4499_), .Y(_4503_) );
OAI21X1 OAI21X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_4501_), .B(_4502_), .C(_4503_), .Y(_4504_) );
AOI21X1 AOI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_4500_), .B(_4504_), .C(bloque_datos_52_bF_buf3_), .Y(_4505_) );
INVX1 INVX1_1126 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf2_), .Y(_4506_) );
NAND3X1 NAND3X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_4503_), .B(_4490_), .C(_4494_), .Y(_4507_) );
OAI21X1 OAI21X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_4501_), .B(_4502_), .C(_4499_), .Y(_4508_) );
AOI21X1 AOI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_4507_), .B(_4508_), .C(_4506_), .Y(_4509_) );
OAI21X1 OAI21X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_4505_), .B(_4509_), .C(_8202_), .Y(_4510_) );
INVX2 INVX2_281 ( .gnd(gnd), .vdd(vdd), .A(_8202_), .Y(_4511_) );
NAND3X1 NAND3X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_4506_), .B(_4507_), .C(_4508_), .Y(_4512_) );
NAND3X1 NAND3X1_1869 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf1_), .B(_4500_), .C(_4504_), .Y(_4513_) );
NAND3X1 NAND3X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_4511_), .B(_4512_), .C(_4513_), .Y(_4514_) );
NAND3X1 NAND3X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_8200_), .C(_4510_), .Y(_4515_) );
OAI21X1 OAI21X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_8041_), .B(_8037_), .C(_8032_), .Y(_4516_) );
OAI21X1 OAI21X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_4505_), .B(_4509_), .C(_4511_), .Y(_4517_) );
NAND3X1 NAND3X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_8202_), .B(_4512_), .C(_4513_), .Y(_4518_) );
NAND3X1 NAND3X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_4518_), .B(_4517_), .C(_4516_), .Y(_4519_) );
NAND2X1 NAND2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf2_), .B(_4497_), .Y(_4520_) );
OR2X2 OR2X2_180 ( .gnd(gnd), .vdd(vdd), .A(_4497_), .B(bloque_datos_40_bF_buf1_), .Y(_4521_) );
NAND2X1 NAND2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_4520_), .B(_4521_), .Y(_4522_) );
INVX2 INVX2_282 ( .gnd(gnd), .vdd(vdd), .A(_4522_), .Y(_4523_) );
XNOR2X1 XNOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_6425_), .B(_4523_), .Y(_4524_) );
NAND3X1 NAND3X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_4524_), .B(_4515_), .C(_4519_), .Y(_4525_) );
AOI21X1 AOI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_4518_), .B(_4517_), .C(_4516_), .Y(_4526_) );
AOI21X1 AOI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_4510_), .C(_8200_), .Y(_4527_) );
INVX1 INVX1_1127 ( .gnd(gnd), .vdd(vdd), .A(_4524_), .Y(_4528_) );
OAI21X1 OAI21X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_4526_), .B(_4527_), .C(_4528_), .Y(_4529_) );
AOI21X1 AOI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_4525_), .B(_4529_), .C(bloque_datos_68_bF_buf2_), .Y(_4530_) );
INVX1 INVX1_1128 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf1_), .Y(_4531_) );
NAND3X1 NAND3X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_4528_), .B(_4515_), .C(_4519_), .Y(_4532_) );
OAI21X1 OAI21X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_4526_), .B(_4527_), .C(_4524_), .Y(_4533_) );
AOI21X1 AOI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_4532_), .B(_4533_), .C(_4531_), .Y(_4534_) );
OAI21X1 OAI21X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_4530_), .B(_4534_), .C(_8199_), .Y(_4535_) );
NAND3X1 NAND3X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_4531_), .B(_4532_), .C(_4533_), .Y(_4536_) );
NAND3X1 NAND3X1_1877 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf0_), .B(_4525_), .C(_4529_), .Y(_4537_) );
NAND3X1 NAND3X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_8048_), .B(_4536_), .C(_4537_), .Y(_4538_) );
NAND3X1 NAND3X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_8198_), .B(_4538_), .C(_4535_), .Y(_4539_) );
INVX1 INVX1_1129 ( .gnd(gnd), .vdd(vdd), .A(_7966_), .Y(_4540_) );
AOI21X1 AOI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_8043_), .B(_8046_), .C(_7835_), .Y(_4541_) );
OAI21X1 OAI21X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_4541_), .B(_4540_), .C(_8047_), .Y(_4542_) );
OAI21X1 OAI21X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_4530_), .B(_4534_), .C(_8048_), .Y(_4543_) );
NAND3X1 NAND3X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_8199_), .B(_4536_), .C(_4537_), .Y(_4544_) );
NAND3X1 NAND3X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_4542_), .B(_4544_), .C(_4543_), .Y(_4545_) );
NAND2X1 NAND2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf2_), .B(_4522_), .Y(_4546_) );
OR2X2 OR2X2_181 ( .gnd(gnd), .vdd(vdd), .A(_4522_), .B(bloque_datos_56_bF_buf1_), .Y(_4547_) );
NAND2X1 NAND2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_4546_), .B(_4547_), .Y(_4548_) );
INVX2 INVX2_283 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .Y(_4549_) );
XNOR2X1 XNOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_6458_), .B(_4549_), .Y(_4550_) );
NAND3X1 NAND3X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_4550_), .B(_4539_), .C(_4545_), .Y(_4551_) );
AOI21X1 AOI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_4544_), .B(_4543_), .C(_4542_), .Y(_4552_) );
AOI21X1 AOI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_4538_), .B(_4535_), .C(_8198_), .Y(_4553_) );
INVX1 INVX1_1130 ( .gnd(gnd), .vdd(vdd), .A(_4550_), .Y(_4554_) );
OAI21X1 OAI21X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_4552_), .B(_4553_), .C(_4554_), .Y(_4555_) );
AOI21X1 AOI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_4551_), .B(_4555_), .C(bloque_datos_84_bF_buf3_), .Y(_4556_) );
INVX1 INVX1_1131 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf2_), .Y(_4557_) );
NAND3X1 NAND3X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_4554_), .B(_4539_), .C(_4545_), .Y(_4558_) );
OAI21X1 OAI21X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_4552_), .B(_4553_), .C(_4550_), .Y(_4559_) );
AOI21X1 AOI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_4558_), .B(_4559_), .C(_4557_), .Y(_4560_) );
OAI21X1 OAI21X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_4556_), .B(_4560_), .C(_8196_), .Y(_4561_) );
NAND3X1 NAND3X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_4557_), .B(_4558_), .C(_4559_), .Y(_4562_) );
NAND3X1 NAND3X1_1885 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf1_), .B(_4551_), .C(_4555_), .Y(_4563_) );
NAND3X1 NAND3X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_8060_), .B(_4562_), .C(_4563_), .Y(_4564_) );
NAND3X1 NAND3X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_4561_), .B(_4564_), .C(_8195_), .Y(_4565_) );
NAND2X1 NAND2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_8058_), .B(_8064_), .Y(_4566_) );
OAI21X1 OAI21X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_4556_), .B(_4560_), .C(_8060_), .Y(_4567_) );
NAND3X1 NAND3X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_8196_), .B(_4562_), .C(_4563_), .Y(_4568_) );
NAND3X1 NAND3X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_4566_), .B(_4568_), .C(_4567_), .Y(_4569_) );
NOR2X1 NOR2X1_613 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf3_), .B(_4549_), .Y(_4570_) );
NAND2X1 NAND2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf2_), .B(_4549_), .Y(_4571_) );
INVX1 INVX1_1132 ( .gnd(gnd), .vdd(vdd), .A(_4571_), .Y(_4572_) );
NOR2X1 NOR2X1_614 ( .gnd(gnd), .vdd(vdd), .A(_4570_), .B(_4572_), .Y(_4573_) );
XOR2X1 XOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_6491_), .B(_4573_), .Y(_4574_) );
NAND3X1 NAND3X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_4574_), .B(_4569_), .C(_4565_), .Y(_4575_) );
AOI21X1 AOI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_4568_), .B(_4567_), .C(_4566_), .Y(_4576_) );
AOI21X1 AOI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_4564_), .B(_4561_), .C(_8195_), .Y(_4577_) );
INVX1 INVX1_1133 ( .gnd(gnd), .vdd(vdd), .A(_4574_), .Y(_4578_) );
OAI21X1 OAI21X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_4576_), .B(_4577_), .C(_4578_), .Y(_4579_) );
AOI21X1 AOI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_4575_), .B(_4579_), .C(module_1_W_132_), .Y(_4580_) );
INVX1 INVX1_1134 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_132_), .Y(_4581_) );
NAND3X1 NAND3X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_4578_), .B(_4569_), .C(_4565_), .Y(_4582_) );
OAI21X1 OAI21X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_4576_), .B(_4577_), .C(_4574_), .Y(_4583_) );
AOI21X1 AOI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_4582_), .B(_4583_), .C(_4581_), .Y(_4584_) );
OAI21X1 OAI21X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_4580_), .B(_4584_), .C(_8066_), .Y(_4585_) );
INVX2 INVX2_284 ( .gnd(gnd), .vdd(vdd), .A(_8066_), .Y(_4586_) );
NAND3X1 NAND3X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_4581_), .B(_4582_), .C(_4583_), .Y(_4587_) );
NAND3X1 NAND3X1_1893 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_132_), .B(_4575_), .C(_4579_), .Y(_4588_) );
NAND3X1 NAND3X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_4586_), .B(_4587_), .C(_4588_), .Y(_4589_) );
AOI21X1 AOI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_4589_), .B(_4585_), .C(_8194_), .Y(_4590_) );
AND2X2 AND2X2_177 ( .gnd(gnd), .vdd(vdd), .A(_8073_), .B(_8070_), .Y(_4591_) );
OAI21X1 OAI21X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_4580_), .B(_4584_), .C(_4586_), .Y(_4592_) );
NAND3X1 NAND3X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_8066_), .B(_4587_), .C(_4588_), .Y(_4593_) );
AOI21X1 AOI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_4593_), .B(_4592_), .C(_4591_), .Y(_4594_) );
NAND2X1 NAND2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf1_), .B(_4573_), .Y(_4595_) );
OR2X2 OR2X2_182 ( .gnd(gnd), .vdd(vdd), .A(_4573_), .B(bloque_datos_88_bF_buf0_), .Y(_4596_) );
NAND2X1 NAND2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_4595_), .B(_4596_), .Y(_4597_) );
OAI21X1 OAI21X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_4590_), .B(_4594_), .C(_4597_), .Y(_4598_) );
AOI21X1 AOI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_4587_), .B(_4588_), .C(_4586_), .Y(_4599_) );
NOR3X1 NOR3X1_237 ( .gnd(gnd), .vdd(vdd), .A(_4580_), .B(_8066_), .C(_4584_), .Y(_4600_) );
OAI21X1 OAI21X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_4600_), .B(_4599_), .C(_4591_), .Y(_4601_) );
NAND3X1 NAND3X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_8194_), .B(_4589_), .C(_4585_), .Y(_4602_) );
INVX2 INVX2_285 ( .gnd(gnd), .vdd(vdd), .A(_4597_), .Y(_4603_) );
NAND3X1 NAND3X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_4602_), .B(_4603_), .C(_4601_), .Y(_4604_) );
NAND2X1 NAND2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_4598_), .B(_4604_), .Y(_4605_) );
NAND3X1 NAND3X1_1898 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_148_), .B(_6524_), .C(_4605_), .Y(_4606_) );
INVX1 INVX1_1135 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_148_), .Y(_4607_) );
AOI21X1 AOI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_4602_), .B(_4601_), .C(_4597_), .Y(_4608_) );
NAND2X1 NAND2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_4602_), .B(_4601_), .Y(_4609_) );
OAI21X1 OAI21X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_4609_), .B(_4603_), .C(_6524_), .Y(_4610_) );
OAI21X1 OAI21X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_4610_), .B(_4608_), .C(_4607_), .Y(_4611_) );
AOI21X1 AOI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_4606_), .B(_4611_), .C(_8079_), .Y(_4612_) );
OAI21X1 OAI21X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_4610_), .B(_4608_), .C(module_1_W_148_), .Y(_4613_) );
NAND3X1 NAND3X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_4607_), .B(_6524_), .C(_4605_), .Y(_4614_) );
AOI21X1 AOI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_4614_), .B(_4613_), .C(_8078_), .Y(_4615_) );
OAI21X1 OAI21X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_4615_), .B(_4612_), .C(_8193_), .Y(_4616_) );
NAND2X1 NAND2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_8080_), .B(_8084_), .Y(_4617_) );
NAND3X1 NAND3X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_8078_), .B(_4614_), .C(_4613_), .Y(_4618_) );
NAND3X1 NAND3X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_8079_), .B(_4606_), .C(_4611_), .Y(_4619_) );
NAND3X1 NAND3X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_4617_), .B(_4618_), .C(_4619_), .Y(_4620_) );
NAND2X1 NAND2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_136_), .B(_4597_), .Y(_4621_) );
OR2X2 OR2X2_183 ( .gnd(gnd), .vdd(vdd), .A(_4597_), .B(module_1_W_136_), .Y(_4622_) );
NAND2X1 NAND2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_4621_), .B(_4622_), .Y(_4623_) );
NAND3X1 NAND3X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_4620_), .B(_4623_), .C(_4616_), .Y(_4624_) );
NAND2X1 NAND2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_4620_), .B(_4616_), .Y(_4625_) );
INVX2 INVX2_286 ( .gnd(gnd), .vdd(vdd), .A(_4623_), .Y(_4626_) );
AOI21X1 AOI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_4626_), .B(_4625_), .C(_6809_), .Y(_4627_) );
NAND3X1 NAND3X1_1904 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_164_), .B(_4624_), .C(_4627_), .Y(_4628_) );
INVX1 INVX1_1136 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_164_), .Y(_4629_) );
AOI21X1 AOI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_4618_), .B(_4619_), .C(_4617_), .Y(_4630_) );
NAND3X1 NAND3X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_8078_), .B(_4606_), .C(_4611_), .Y(_4631_) );
NAND3X1 NAND3X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_8079_), .B(_4614_), .C(_4613_), .Y(_4632_) );
AOI21X1 AOI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_4631_), .B(_4632_), .C(_8193_), .Y(_4633_) );
OAI21X1 OAI21X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_4630_), .B(_4633_), .C(_4626_), .Y(_4634_) );
NAND3X1 NAND3X1_1907 ( .gnd(gnd), .vdd(vdd), .A(_6557_), .B(_4624_), .C(_4634_), .Y(_4635_) );
NAND2X1 NAND2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_4629_), .B(_4635_), .Y(_4636_) );
AOI21X1 AOI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_4636_), .B(_4628_), .C(_8089_), .Y(_4637_) );
INVX1 INVX1_1137 ( .gnd(gnd), .vdd(vdd), .A(_8089_), .Y(_4638_) );
NAND2X1 NAND2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_164_), .B(_4635_), .Y(_4639_) );
NAND3X1 NAND3X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_4629_), .B(_4624_), .C(_4627_), .Y(_4640_) );
AOI21X1 AOI21X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_4639_), .B(_4640_), .C(_4638_), .Y(_4641_) );
OAI21X1 OAI21X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_4641_), .B(_4637_), .C(_8192_), .Y(_4642_) );
NAND3X1 NAND3X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_4638_), .B(_4639_), .C(_4640_), .Y(_4643_) );
NAND3X1 NAND3X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_8089_), .B(_4636_), .C(_4628_), .Y(_4644_) );
NAND3X1 NAND3X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_8191_), .B(_4643_), .C(_4644_), .Y(_4645_) );
NAND2X1 NAND2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_152_), .B(_4623_), .Y(_4646_) );
OR2X2 OR2X2_184 ( .gnd(gnd), .vdd(vdd), .A(_4623_), .B(module_1_W_152_), .Y(_4647_) );
NAND2X1 NAND2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_4646_), .B(_4647_), .Y(_4648_) );
NAND3X1 NAND3X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_4645_), .B(_4648_), .C(_4642_), .Y(_4649_) );
AOI21X1 AOI21X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_4645_), .B(_4642_), .C(_4648_), .Y(_4650_) );
NOR2X1 NOR2X1_615 ( .gnd(gnd), .vdd(vdd), .A(_6787_), .B(_4650_), .Y(_4651_) );
NAND3X1 NAND3X1_1913 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_180_), .B(_4649_), .C(_4651_), .Y(_4652_) );
INVX1 INVX1_1138 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_180_), .Y(_4653_) );
NAND2X1 NAND2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_6590_), .B(_4649_), .Y(_4654_) );
OAI21X1 OAI21X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_4654_), .B(_4650_), .C(_4653_), .Y(_4655_) );
AOI21X1 AOI21X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_4655_), .B(_4652_), .C(_8102_), .Y(_4656_) );
OAI21X1 OAI21X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_4654_), .B(_4650_), .C(module_1_W_180_), .Y(_4657_) );
NAND3X1 NAND3X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_4653_), .B(_4649_), .C(_4651_), .Y(_4658_) );
AOI21X1 AOI21X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_4657_), .B(_4658_), .C(_8101_), .Y(_4659_) );
OAI21X1 OAI21X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_4659_), .B(_4656_), .C(_8189_), .Y(_4660_) );
OAI21X1 OAI21X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_8109_), .B(_7956_), .C(_8103_), .Y(_4661_) );
NAND3X1 NAND3X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_8101_), .B(_4657_), .C(_4658_), .Y(_4662_) );
NAND3X1 NAND3X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_8102_), .B(_4655_), .C(_4652_), .Y(_4663_) );
NAND3X1 NAND3X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_4662_), .B(_4661_), .C(_4663_), .Y(_4664_) );
NAND2X1 NAND2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_168_), .B(_4648_), .Y(_4665_) );
OR2X2 OR2X2_185 ( .gnd(gnd), .vdd(vdd), .A(_4648_), .B(module_1_W_168_), .Y(_4666_) );
NAND2X1 NAND2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_4665_), .B(_4666_), .Y(_4667_) );
NAND3X1 NAND3X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_4664_), .B(_4667_), .C(_4660_), .Y(_4668_) );
NAND2X1 NAND2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_4664_), .B(_4660_), .Y(_4669_) );
INVX2 INVX2_287 ( .gnd(gnd), .vdd(vdd), .A(_4667_), .Y(_4670_) );
AOI21X1 AOI21X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_4670_), .B(_4669_), .C(_6754_), .Y(_4671_) );
NAND3X1 NAND3X1_1919 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_196_), .B(_4668_), .C(_4671_), .Y(_4672_) );
INVX1 INVX1_1139 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_196_), .Y(_4673_) );
AOI21X1 AOI21X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_4662_), .B(_4663_), .C(_4661_), .Y(_4674_) );
NOR3X1 NOR3X1_238 ( .gnd(gnd), .vdd(vdd), .A(_4656_), .B(_8189_), .C(_4659_), .Y(_4675_) );
OAI21X1 OAI21X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_4675_), .B(_4674_), .C(_4670_), .Y(_4676_) );
NAND3X1 NAND3X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_6623_), .B(_4668_), .C(_4676_), .Y(_4677_) );
NAND2X1 NAND2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_4673_), .B(_4677_), .Y(_4678_) );
AOI21X1 AOI21X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_4672_), .B(_4678_), .C(_8114_), .Y(_4679_) );
INVX1 INVX1_1140 ( .gnd(gnd), .vdd(vdd), .A(_8107_), .Y(_4680_) );
NAND2X1 NAND2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_8110_), .B(_4680_), .Y(_4681_) );
NOR2X1 NOR2X1_616 ( .gnd(gnd), .vdd(vdd), .A(_7955_), .B(_4681_), .Y(_4682_) );
NAND2X1 NAND2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_196_), .B(_4677_), .Y(_4683_) );
NAND3X1 NAND3X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_4673_), .B(_4668_), .C(_4671_), .Y(_4684_) );
AOI21X1 AOI21X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_4684_), .B(_4683_), .C(_4682_), .Y(_4685_) );
OAI21X1 OAI21X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_4679_), .B(_4685_), .C(_8187_), .Y(_4686_) );
OAI21X1 OAI21X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .B(_7953_), .C(_8116_), .Y(_4687_) );
NAND3X1 NAND3X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_4682_), .B(_4684_), .C(_4683_), .Y(_4688_) );
NAND3X1 NAND3X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_8114_), .B(_4672_), .C(_4678_), .Y(_4689_) );
NAND3X1 NAND3X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_4688_), .B(_4689_), .C(_4687_), .Y(_4690_) );
NAND2X1 NAND2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_4690_), .B(_4686_), .Y(_4691_) );
NAND2X1 NAND2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_184_), .B(_4667_), .Y(_4692_) );
OR2X2 OR2X2_186 ( .gnd(gnd), .vdd(vdd), .A(_4667_), .B(module_1_W_184_), .Y(_4693_) );
NAND2X1 NAND2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_4692_), .B(_4693_), .Y(_4694_) );
INVX2 INVX2_288 ( .gnd(gnd), .vdd(vdd), .A(_4694_), .Y(_4695_) );
OR2X2 OR2X2_187 ( .gnd(gnd), .vdd(vdd), .A(_4691_), .B(_4695_), .Y(_4696_) );
AOI21X1 AOI21X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_4690_), .B(_4686_), .C(_4694_), .Y(_4697_) );
NOR2X1 NOR2X1_617 ( .gnd(gnd), .vdd(vdd), .A(_6733_), .B(_4697_), .Y(_4698_) );
NAND3X1 NAND3X1_1925 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_212_), .B(_4696_), .C(_4698_), .Y(_4699_) );
INVX1 INVX1_1141 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_212_), .Y(_4700_) );
OAI21X1 OAI21X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_4691_), .B(_4695_), .C(_6656_), .Y(_4701_) );
OAI21X1 OAI21X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_4701_), .B(_4697_), .C(_4700_), .Y(_4702_) );
AOI21X1 AOI21X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_4702_), .B(_4699_), .C(_8132_), .Y(_4703_) );
OAI21X1 OAI21X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_4701_), .B(_4697_), .C(module_1_W_212_), .Y(_4704_) );
NAND3X1 NAND3X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_4700_), .B(_4696_), .C(_4698_), .Y(_4705_) );
AOI21X1 AOI21X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_4704_), .B(_4705_), .C(_8129_), .Y(_4706_) );
OAI21X1 OAI21X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_4703_), .B(_4706_), .C(_8185_), .Y(_4707_) );
NAND3X1 NAND3X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_7910_), .B(_8124_), .C(_8132_), .Y(_4708_) );
OAI21X1 OAI21X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_8136_), .B(_8133_), .C(_4708_), .Y(_4709_) );
NAND3X1 NAND3X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_8129_), .B(_4704_), .C(_4705_), .Y(_4710_) );
NAND3X1 NAND3X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_8132_), .B(_4702_), .C(_4699_), .Y(_4711_) );
INVX1 INVX1_1142 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_0_), .Y(_8467_) );
INVX4 INVX4_7 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf2), .Y(_8468_) );
NAND2X1 NAND2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(nonce_iniciales[32]), .B(_8468_), .Y(_8288_) );
OAI21X1 OAI21X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_8467_), .B(_8468_), .C(_8288_), .Y(_8287__0_) );
INVX1 INVX1_1143 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_1_), .Y(_8289_) );
NAND2X1 NAND2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(nonce_iniciales[33]), .B(_8468_), .Y(_8290_) );
OAI21X1 OAI21X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_8468_), .B(_8289_), .C(_8290_), .Y(_8287__1_) );
NAND2X1 NAND2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_5_), .B(module_1_W_4_), .Y(_8291_) );
NAND2X1 NAND2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_7_), .B(module_1_W_6_), .Y(_8292_) );
NOR2X1 NOR2X1_618 ( .gnd(gnd), .vdd(vdd), .A(_8291_), .B(_8292_), .Y(_8293_) );
NAND2X1 NAND2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_25_), .B(module_1_W_24_), .Y(_8294_) );
NAND2X1 NAND2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_27_), .B(module_1_W_26_), .Y(_8295_) );
NOR2X1 NOR2X1_619 ( .gnd(gnd), .vdd(vdd), .A(_8294_), .B(_8295_), .Y(_8296_) );
INVX1 INVX1_1144 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_2_), .Y(_8297_) );
OAI21X1 OAI21X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_8467_), .B(_8289_), .C(_8297_), .Y(_8298_) );
NAND3X1 NAND3X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_8298_), .B(_8293_), .C(_8296_), .Y(_8299_) );
INVX1 INVX1_1145 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_29_), .Y(_8300_) );
INVX1 INVX1_1146 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_28_), .Y(_8301_) );
NOR2X1 NOR2X1_620 ( .gnd(gnd), .vdd(vdd), .A(_8300_), .B(_8301_), .Y(_8302_) );
INVX1 INVX1_1147 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_31_), .Y(_8303_) );
INVX1 INVX1_1148 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_30_), .Y(_8304_) );
NOR2X1 NOR2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_8303_), .B(_8304_), .Y(_8305_) );
NAND3X1 NAND3X1_1931 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_3_), .B(_8302_), .C(_8305_), .Y(_8306_) );
NOR2X1 NOR2X1_622 ( .gnd(gnd), .vdd(vdd), .A(_8306_), .B(_8299_), .Y(_8307_) );
NAND2X1 NAND2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_17_), .B(module_1_W_16_), .Y(_8308_) );
NAND2X1 NAND2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_19_), .B(module_1_W_18_), .Y(_8309_) );
NOR2X1 NOR2X1_623 ( .gnd(gnd), .vdd(vdd), .A(_8308_), .B(_8309_), .Y(_8310_) );
NAND2X1 NAND2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_22_), .B(module_1_W_21_), .Y(_8311_) );
NAND2X1 NAND2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_23_), .B(module_1_W_20_), .Y(_8312_) );
NOR2X1 NOR2X1_624 ( .gnd(gnd), .vdd(vdd), .A(_8311_), .B(_8312_), .Y(_8313_) );
NAND2X1 NAND2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_8310_), .B(_8313_), .Y(_8314_) );
NAND2X1 NAND2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_9_), .B(module_1_W_8_), .Y(_8315_) );
NAND2X1 NAND2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_11_), .B(module_1_W_10_), .Y(_8316_) );
NOR2X1 NOR2X1_625 ( .gnd(gnd), .vdd(vdd), .A(_8315_), .B(_8316_), .Y(_8317_) );
NAND2X1 NAND2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_15_), .B(module_1_W_14_), .Y(_8318_) );
NAND2X1 NAND2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_13_), .B(module_1_W_12_), .Y(_8319_) );
NOR2X1 NOR2X1_626 ( .gnd(gnd), .vdd(vdd), .A(_8318_), .B(_8319_), .Y(_8320_) );
NAND2X1 NAND2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_8317_), .B(_8320_), .Y(_8321_) );
NOR2X1 NOR2X1_627 ( .gnd(gnd), .vdd(vdd), .A(_8314_), .B(_8321_), .Y(_8322_) );
AOI21X1 AOI21X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_8322_), .B(_8307_), .C(_8468_), .Y(_8323_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_2_), .B(nonce_iniciales[34]), .S(inicio_bF_buf3), .Y(_8324_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_2_), .B(_8324_), .S(_8323__bF_buf2), .Y(_8287__2_) );
NAND2X1 NAND2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_2_), .B(module_1_W_3_), .Y(_8325_) );
INVX1 INVX1_1149 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_3_), .Y(_8326_) );
NAND2X1 NAND2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_8297_), .B(_8326_), .Y(_8327_) );
NAND2X1 NAND2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_8325_), .B(_8327_), .Y(_8328_) );
NOR2X1 NOR2X1_628 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf2), .B(nonce_iniciales[35]), .Y(_8329_) );
AOI21X1 AOI21X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_8328_), .B(_8323__bF_buf2), .C(_8329_), .Y(_8287__3_) );
XOR2X1 XOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_8325_), .B(module_1_W_4_), .Y(_8330_) );
NOR2X1 NOR2X1_629 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf2), .B(nonce_iniciales[36]), .Y(_8331_) );
AOI21X1 AOI21X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_8330_), .B(_8323__bF_buf3), .C(_8331_), .Y(_8287__4_) );
AND2X2 AND2X2_178 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_2_), .B(module_1_W_3_), .Y(_8332_) );
NAND2X1 NAND2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_4_), .B(_8332_), .Y(_8333_) );
XOR2X1 XOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_8333_), .B(module_1_W_5_), .Y(_8334_) );
NOR2X1 NOR2X1_630 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf2), .B(nonce_iniciales[37]), .Y(_8335_) );
AOI21X1 AOI21X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_8334_), .B(_8323__bF_buf3), .C(_8335_), .Y(_8287__5_) );
NOR2X1 NOR2X1_631 ( .gnd(gnd), .vdd(vdd), .A(_8291_), .B(_8325_), .Y(_8336_) );
XNOR2X1 XNOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_8336_), .B(module_1_W_6_), .Y(_8337_) );
NOR2X1 NOR2X1_632 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf3), .B(nonce_iniciales[38]), .Y(_8338_) );
AOI21X1 AOI21X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_8337_), .B(_8323__bF_buf2), .C(_8338_), .Y(_8287__6_) );
NOR2X1 NOR2X1_633 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf3), .B(nonce_iniciales[39]), .Y(_8339_) );
NAND2X1 NAND2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_6_), .B(_8336_), .Y(_8340_) );
XOR2X1 XOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_8340_), .B(module_1_W_7_), .Y(_8341_) );
AOI21X1 AOI21X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_8341_), .B(_8323__bF_buf3), .C(_8339_), .Y(_8287__7_) );
NOR3X1 NOR3X1_239 ( .gnd(gnd), .vdd(vdd), .A(_8291_), .B(_8292_), .C(_8325_), .Y(_8342_) );
XNOR2X1 XNOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_8342_), .B(module_1_W_8_), .Y(_8343_) );
NOR2X1 NOR2X1_634 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf2), .B(nonce_iniciales[40]), .Y(_8344_) );
AOI21X1 AOI21X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_8343_), .B(_8323__bF_buf2), .C(_8344_), .Y(_8287__8_) );
AND2X2 AND2X2_179 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_5_), .B(module_1_W_4_), .Y(_8345_) );
AND2X2 AND2X2_180 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_7_), .B(module_1_W_6_), .Y(_8346_) );
NAND3X1 NAND3X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_8345_), .B(_8346_), .C(_8332_), .Y(_8347_) );
INVX1 INVX1_1150 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_9_), .Y(_8348_) );
INVX1 INVX1_1151 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_8_), .Y(_8349_) );
OAI21X1 OAI21X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_8347_), .B(_8349_), .C(_8348_), .Y(_8350_) );
OAI21X1 OAI21X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_8315_), .B(_8347_), .C(_8350_), .Y(_8351_) );
NOR2X1 NOR2X1_635 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf2), .B(nonce_iniciales[41]), .Y(_8352_) );
AOI21X1 AOI21X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_8351_), .B(_8323__bF_buf3), .C(_8352_), .Y(_8287__9_) );
NOR2X1 NOR2X1_636 ( .gnd(gnd), .vdd(vdd), .A(_8315_), .B(_8347_), .Y(_8353_) );
XNOR2X1 XNOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_8353_), .B(module_1_W_10_), .Y(_8354_) );
NOR2X1 NOR2X1_637 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf2), .B(nonce_iniciales[42]), .Y(_8355_) );
AOI21X1 AOI21X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_8354_), .B(_8323__bF_buf2), .C(_8355_), .Y(_8287__10_) );
NOR2X1 NOR2X1_638 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[43]), .Y(_8356_) );
NAND2X1 NAND2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_10_), .B(_8353_), .Y(_8357_) );
OR2X2 OR2X2_188 ( .gnd(gnd), .vdd(vdd), .A(_8357_), .B(module_1_W_11_), .Y(_8358_) );
NAND2X1 NAND2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_8322_), .B(_8307_), .Y(_8359_) );
NAND2X1 NAND2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf2), .B(_8359_), .Y(_8360_) );
AOI21X1 AOI21X1_1187 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_11_), .B(_8357_), .C(_8360_), .Y(_8361_) );
AOI21X1 AOI21X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_8358_), .B(_8361_), .C(_8356_), .Y(_8287__11_) );
INVX2 INVX2_289 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_12_), .Y(_8362_) );
NAND2X1 NAND2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_8317_), .B(_8342_), .Y(_8363_) );
XNOR2X1 XNOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_8363_), .B(_8362_), .Y(_8364_) );
NOR2X1 NOR2X1_639 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[44]), .Y(_8365_) );
AOI21X1 AOI21X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_8364_), .B(_8323__bF_buf1), .C(_8365_), .Y(_8287__12_) );
NOR2X1 NOR2X1_640 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[45]), .Y(_8366_) );
INVX1 INVX1_1152 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_13_), .Y(_8367_) );
NAND3X1 NAND3X1_1933 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_11_), .B(module_1_W_10_), .C(_8353_), .Y(_8368_) );
NOR2X1 NOR2X1_641 ( .gnd(gnd), .vdd(vdd), .A(_8362_), .B(_8368_), .Y(_8369_) );
NAND2X1 NAND2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_8367_), .B(_8369_), .Y(_8370_) );
OAI21X1 OAI21X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_8363_), .B(_8362_), .C(module_1_W_13_), .Y(_8371_) );
AND2X2 AND2X2_181 ( .gnd(gnd), .vdd(vdd), .A(_8323__bF_buf0), .B(_8371_), .Y(_8372_) );
AOI21X1 AOI21X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_8370_), .B(_8372_), .C(_8366_), .Y(_8287__13_) );
INVX2 INVX2_290 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_14_), .Y(_8373_) );
OR2X2 OR2X2_189 ( .gnd(gnd), .vdd(vdd), .A(_8363_), .B(_8319_), .Y(_8374_) );
XNOR2X1 XNOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_8374_), .B(_8373_), .Y(_8375_) );
NOR2X1 NOR2X1_642 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[46]), .Y(_8376_) );
AOI21X1 AOI21X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_8323__bF_buf0), .B(_8375_), .C(_8376_), .Y(_8287__14_) );
NOR2X1 NOR2X1_643 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[47]), .Y(_8377_) );
INVX1 INVX1_1153 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_15_), .Y(_8378_) );
NOR2X1 NOR2X1_644 ( .gnd(gnd), .vdd(vdd), .A(_8319_), .B(_8368_), .Y(_8379_) );
NAND3X1 NAND3X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_8378_), .B(module_1_W_14_), .C(_8379_), .Y(_8380_) );
OAI21X1 OAI21X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_8374_), .B(_8373_), .C(module_1_W_15_), .Y(_8381_) );
AND2X2 AND2X2_182 ( .gnd(gnd), .vdd(vdd), .A(_8381_), .B(_8323__bF_buf2), .Y(_8382_) );
AOI21X1 AOI21X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_8380_), .B(_8382_), .C(_8377_), .Y(_8287__15_) );
OR2X2 OR2X2_190 ( .gnd(gnd), .vdd(vdd), .A(_8315_), .B(_8316_), .Y(_8383_) );
OR2X2 OR2X2_191 ( .gnd(gnd), .vdd(vdd), .A(_8318_), .B(_8319_), .Y(_8384_) );
NOR3X1 NOR3X1_240 ( .gnd(gnd), .vdd(vdd), .A(_8384_), .B(_8383_), .C(_8347_), .Y(_8385_) );
NAND2X1 NAND2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_16_), .B(_8385_), .Y(_8386_) );
INVX1 INVX1_1154 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_16_), .Y(_8387_) );
OAI21X1 OAI21X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_8321_), .B(_8347_), .C(_8387_), .Y(_8388_) );
NAND2X1 NAND2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_8388_), .B(_8386_), .Y(_8389_) );
NOR2X1 NOR2X1_645 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[48]), .Y(_8390_) );
AOI21X1 AOI21X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_8323__bF_buf1), .B(_8389_), .C(_8390_), .Y(_8287__16_) );
NAND3X1 NAND3X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_8317_), .B(_8320_), .C(_8342_), .Y(_8391_) );
NOR2X1 NOR2X1_646 ( .gnd(gnd), .vdd(vdd), .A(_8387_), .B(_8391_), .Y(_8392_) );
XNOR2X1 XNOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_8392_), .B(module_1_W_17_), .Y(_8393_) );
NOR2X1 NOR2X1_647 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[49]), .Y(_8394_) );
AOI21X1 AOI21X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_8323__bF_buf1), .B(_8393_), .C(_8394_), .Y(_8287__17_) );
INVX1 INVX1_1155 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_18_), .Y(_8395_) );
INVX1 INVX1_1156 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_17_), .Y(_8396_) );
OAI21X1 OAI21X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_8386_), .B(_8396_), .C(_8395_), .Y(_8397_) );
NAND3X1 NAND3X1_1936 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_18_), .B(module_1_W_17_), .C(_8392_), .Y(_8398_) );
NAND2X1 NAND2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_8398_), .B(_8397_), .Y(_8399_) );
NOR2X1 NOR2X1_648 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[50]), .Y(_8400_) );
AOI21X1 AOI21X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_8323__bF_buf1), .B(_8399_), .C(_8400_), .Y(_8287__18_) );
NOR2X1 NOR2X1_649 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[51]), .Y(_8401_) );
OR2X2 OR2X2_192 ( .gnd(gnd), .vdd(vdd), .A(_8398_), .B(module_1_W_19_), .Y(_8402_) );
AOI21X1 AOI21X1_1196 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_19_), .B(_8398_), .C(_8360_), .Y(_8403_) );
AOI21X1 AOI21X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_8402_), .B(_8403_), .C(_8401_), .Y(_8287__19_) );
INVX1 INVX1_1157 ( .gnd(gnd), .vdd(vdd), .A(_8310_), .Y(_8404_) );
NOR2X1 NOR2X1_650 ( .gnd(gnd), .vdd(vdd), .A(_8404_), .B(_8391_), .Y(_8405_) );
NAND2X1 NAND2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_20_), .B(_8405_), .Y(_8406_) );
INVX2 INVX2_291 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_20_), .Y(_8407_) );
OAI21X1 OAI21X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_8391_), .B(_8404_), .C(_8407_), .Y(_8408_) );
NAND2X1 NAND2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_8408_), .B(_8406_), .Y(_8409_) );
NOR2X1 NOR2X1_651 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf2), .B(nonce_iniciales[52]), .Y(_8410_) );
AOI21X1 AOI21X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_8323__bF_buf3), .B(_8409_), .C(_8410_), .Y(_8287__20_) );
INVX1 INVX1_1158 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_21_), .Y(_8411_) );
INVX1 INVX1_1159 ( .gnd(gnd), .vdd(vdd), .A(_8359_), .Y(_8412_) );
NAND2X1 NAND2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_8310_), .B(_8385_), .Y(_8413_) );
NOR2X1 NOR2X1_652 ( .gnd(gnd), .vdd(vdd), .A(_8407_), .B(_8413_), .Y(_8414_) );
AOI21X1 AOI21X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_8411_), .B(_8414_), .C(_8412_), .Y(_8415_) );
AOI21X1 AOI21X1_1200 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_21_), .B(_8406_), .C(_8468_), .Y(_8416_) );
NOR2X1 NOR2X1_653 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[53]), .Y(_8417_) );
AOI21X1 AOI21X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_8416_), .B(_8415_), .C(_8417_), .Y(_8287__21_) );
NOR2X1 NOR2X1_654 ( .gnd(gnd), .vdd(vdd), .A(_8411_), .B(_8407_), .Y(_8418_) );
INVX1 INVX1_1160 ( .gnd(gnd), .vdd(vdd), .A(_8418_), .Y(_8419_) );
OAI21X1 OAI21X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_8413_), .B(_8419_), .C(module_1_W_22_), .Y(_8420_) );
INVX1 INVX1_1161 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_22_), .Y(_8421_) );
NAND3X1 NAND3X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_8421_), .B(_8418_), .C(_8405_), .Y(_8422_) );
AND2X2 AND2X2_183 ( .gnd(gnd), .vdd(vdd), .A(_8420_), .B(_8422_), .Y(_8423_) );
NOR2X1 NOR2X1_655 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf2), .B(nonce_iniciales[54]), .Y(_8424_) );
AOI21X1 AOI21X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_8323__bF_buf3), .B(_8423_), .C(_8424_), .Y(_8287__22_) );
NOR2X1 NOR2X1_656 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf2), .B(nonce_iniciales[55]), .Y(_8425_) );
INVX1 INVX1_1162 ( .gnd(gnd), .vdd(vdd), .A(_8311_), .Y(_8426_) );
NAND3X1 NAND3X1_1938 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_20_), .B(_8426_), .C(_8405_), .Y(_8427_) );
OR2X2 OR2X2_193 ( .gnd(gnd), .vdd(vdd), .A(_8427_), .B(module_1_W_23_), .Y(_8428_) );
AOI21X1 AOI21X1_1203 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_23_), .B(_8427_), .C(_8360_), .Y(_8429_) );
AOI21X1 AOI21X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_8428_), .B(_8429_), .C(_8425_), .Y(_8287__23_) );
NOR2X1 NOR2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_8314_), .B(_8391_), .Y(_8430_) );
XNOR2X1 XNOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_8430_), .B(module_1_W_24_), .Y(_8431_) );
NOR2X1 NOR2X1_658 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf6), .B(nonce_iniciales[56]), .Y(_8432_) );
AOI21X1 AOI21X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_8323__bF_buf0), .B(_8431_), .C(_8432_), .Y(_8287__24_) );
INVX1 INVX1_1163 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_25_), .Y(_8433_) );
AND2X2 AND2X2_184 ( .gnd(gnd), .vdd(vdd), .A(_8430_), .B(module_1_W_24_), .Y(_8434_) );
AOI21X1 AOI21X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_8433_), .B(_8434_), .C(_8412_), .Y(_8435_) );
NAND2X1 NAND2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_24_), .B(_8430_), .Y(_8436_) );
AOI21X1 AOI21X1_1207 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_25_), .B(_8436_), .C(_8468_), .Y(_8437_) );
NOR2X1 NOR2X1_659 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf6), .B(nonce_iniciales[57]), .Y(_8438_) );
AOI21X1 AOI21X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_8437_), .B(_8435_), .C(_8438_), .Y(_8287__25_) );
NOR3X1 NOR3X1_241 ( .gnd(gnd), .vdd(vdd), .A(_8294_), .B(_8314_), .C(_8391_), .Y(_8439_) );
XNOR2X1 XNOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_8439_), .B(module_1_W_26_), .Y(_8440_) );
NOR2X1 NOR2X1_660 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf6), .B(nonce_iniciales[58]), .Y(_8441_) );
AOI21X1 AOI21X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_8323__bF_buf0), .B(_8440_), .C(_8441_), .Y(_8287__26_) );
NOR2X1 NOR2X1_661 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf6), .B(nonce_iniciales[59]), .Y(_8442_) );
AND2X2 AND2X2_185 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_26_), .B(module_1_W_25_), .Y(_8443_) );
NAND3X1 NAND3X1_1939 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_24_), .B(_8443_), .C(_8430_), .Y(_8444_) );
OR2X2 OR2X2_194 ( .gnd(gnd), .vdd(vdd), .A(_8444_), .B(module_1_W_27_), .Y(_8445_) );
AOI21X1 AOI21X1_1210 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_27_), .B(_8444_), .C(_8360_), .Y(_8446_) );
AOI21X1 AOI21X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_8445_), .B(_8446_), .C(_8442_), .Y(_8287__27_) );
INVX1 INVX1_1164 ( .gnd(gnd), .vdd(vdd), .A(_8296_), .Y(_8447_) );
NOR3X1 NOR3X1_242 ( .gnd(gnd), .vdd(vdd), .A(_8447_), .B(_8314_), .C(_8391_), .Y(_8448_) );
NAND2X1 NAND2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_28_), .B(_8448_), .Y(_8449_) );
INVX1 INVX1_1165 ( .gnd(gnd), .vdd(vdd), .A(_8314_), .Y(_8450_) );
NAND3X1 NAND3X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_8296_), .B(_8450_), .C(_8385_), .Y(_8451_) );
NAND2X1 NAND2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_8301_), .B(_8451_), .Y(_8452_) );
NAND2X1 NAND2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_8449_), .B(_8452_), .Y(_8453_) );
NOR2X1 NOR2X1_662 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf6), .B(nonce_iniciales[60]), .Y(_8454_) );
AOI21X1 AOI21X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_8323__bF_buf0), .B(_8453_), .C(_8454_), .Y(_8287__28_) );
NOR2X1 NOR2X1_663 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf6), .B(nonce_iniciales[61]), .Y(_8455_) );
OR2X2 OR2X2_195 ( .gnd(gnd), .vdd(vdd), .A(_8449_), .B(module_1_W_29_), .Y(_8456_) );
AOI21X1 AOI21X1_1213 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_29_), .B(_8449_), .C(_8360_), .Y(_8457_) );
AOI21X1 AOI21X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_8456_), .B(_8457_), .C(_8455_), .Y(_8287__29_) );
NAND3X1 NAND3X1_1941 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_30_), .B(_8302_), .C(_8448_), .Y(_8458_) );
INVX1 INVX1_1166 ( .gnd(gnd), .vdd(vdd), .A(_8302_), .Y(_8459_) );
OAI21X1 OAI21X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_8451_), .B(_8459_), .C(_8304_), .Y(_8460_) );
NAND2X1 NAND2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_8458_), .B(_8460_), .Y(_8461_) );
NOR2X1 NOR2X1_664 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[62]), .Y(_8462_) );
AOI21X1 AOI21X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_8323__bF_buf1), .B(_8461_), .C(_8462_), .Y(_8287__30_) );
NOR2X1 NOR2X1_665 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf9), .B(nonce_iniciales[63]), .Y(_8463_) );
NOR2X1 NOR2X1_666 ( .gnd(gnd), .vdd(vdd), .A(_8459_), .B(_8451_), .Y(_8464_) );
NAND3X1 NAND3X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_8303_), .B(module_1_W_30_), .C(_8464_), .Y(_8465_) );
AOI21X1 AOI21X1_1216 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_31_), .B(_8458_), .C(_8360_), .Y(_8466_) );
AOI21X1 AOI21X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_8465_), .B(_8466_), .C(_8463_), .Y(_8287__31_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_8287__0_), .Q(module_1_W_0_) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_8287__1_), .Q(module_1_W_1_) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_8287__2_), .Q(module_1_W_2_) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_8287__3_), .Q(module_1_W_3_) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_8287__4_), .Q(module_1_W_4_) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_8287__5_), .Q(module_1_W_5_) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_8287__6_), .Q(module_1_W_6_) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_8287__7_), .Q(module_1_W_7_) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_8287__8_), .Q(module_1_W_8_) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_8287__9_), .Q(module_1_W_9_) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_8287__10_), .Q(module_1_W_10_) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8287__11_), .Q(module_1_W_11_) );
DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8287__12_), .Q(module_1_W_12_) );
DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8287__13_), .Q(module_1_W_13_) );
DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8287__14_), .Q(module_1_W_14_) );
DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8287__15_), .Q(module_1_W_15_) );
DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8287__16_), .Q(module_1_W_16_) );
DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8287__17_), .Q(module_1_W_17_) );
DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8287__18_), .Q(module_1_W_18_) );
DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8287__19_), .Q(module_1_W_19_) );
DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_8287__20_), .Q(module_1_W_20_) );
DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_8287__21_), .Q(module_1_W_21_) );
DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_8287__22_), .Q(module_1_W_22_) );
DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_8287__23_), .Q(module_1_W_23_) );
DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_8287__24_), .Q(module_1_W_24_) );
DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8287__25_), .Q(module_1_W_25_) );
DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_8287__26_), .Q(module_1_W_26_) );
DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_8287__27_), .Q(module_1_W_27_) );
DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_8287__28_), .Q(module_1_W_28_) );
DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_8287__29_), .Q(module_1_W_29_) );
DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8287__30_), .Q(module_1_W_30_) );
DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_8287__31_), .Q(module_1_W_31_) );
INVX1 INVX1_1167 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_8506_) );
INVX1 INVX1_1168 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .Y(_8507_) );
INVX1 INVX1_1169 ( .gnd(gnd), .vdd(vdd), .A(target[0]), .Y(_8508_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_8507_), .B(gnd), .C(_8508_), .D(vdd), .Y(_8509_) );
OAI21X1 OAI21X1_1360 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .B(_8506_), .C(_8509_), .Y(_8510_) );
XOR2X1 XOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(vdd), .Y(_8511_) );
INVX2 INVX2_292 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .Y(_8512_) );
INVX1 INVX1_1170 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_8513_) );
NAND2X1 NAND2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_8512_), .B(_8513_), .Y(_8514_) );
NAND2X1 NAND2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(gnd), .Y(_8515_) );
AOI21X1 AOI21X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_8514_), .B(_8515_), .C(_8511_), .Y(_8516_) );
INVX1 INVX1_1171 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .Y(_8517_) );
NAND2X1 NAND2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_8517_), .Y(_8518_) );
NAND2X1 NAND2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_8512_), .Y(_8519_) );
OAI21X1 OAI21X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_8511_), .B(_8519_), .C(_8518_), .Y(_8520_) );
AOI21X1 AOI21X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_8510_), .B(_8516_), .C(_8520_), .Y(_8521_) );
INVX1 INVX1_1172 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_15_), .Y(_8522_) );
INVX1 INVX1_1173 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_14_), .Y(_8523_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_8522_), .B(target[7]), .C(target[6]), .D(_8523_), .Y(_8524_) );
INVX4 INVX4_8 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .Y(_8525_) );
INVX2 INVX2_293 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .Y(_8526_) );
OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_8525_), .B(module_1_H_15_), .C(_8526_), .D(module_1_H_14_), .Y(_8527_) );
NOR2X1 NOR2X1_667 ( .gnd(gnd), .vdd(vdd), .A(_8524_), .B(_8527_), .Y(_8528_) );
INVX2 INVX2_294 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_13_), .Y(_8529_) );
INVX1 INVX1_1174 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_12_), .Y(_8530_) );
OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_8529_), .B(target[5]), .C(target[4]), .D(_8530_), .Y(_8531_) );
INVX2 INVX2_295 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .Y(_8532_) );
INVX1 INVX1_1175 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .Y(_8533_) );
OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_8532_), .B(module_1_H_13_), .C(_8533_), .D(module_1_H_12_), .Y(_8534_) );
NOR2X1 NOR2X1_668 ( .gnd(gnd), .vdd(vdd), .A(_8531_), .B(_8534_), .Y(_8535_) );
NAND2X1 NAND2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_8528_), .B(_8535_), .Y(_8536_) );
NAND2X1 NAND2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .B(_8529_), .Y(_8537_) );
NAND3X1 NAND3X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_8531_), .B(_8537_), .C(_8528_), .Y(_8538_) );
OAI21X1 OAI21X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_8521_), .B(_8536_), .C(_8538_), .Y(_8539_) );
INVX1 INVX1_1176 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_17_), .Y(_8540_) );
OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_8507_), .B(module_1_H_17_), .C(_8508_), .D(module_1_H_16_), .Y(_8541_) );
OAI21X1 OAI21X1_1363 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .B(_8540_), .C(_8541_), .Y(_8542_) );
XOR2X1 XOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(module_1_H_19_), .Y(_8543_) );
INVX1 INVX1_1177 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_18_), .Y(_8544_) );
NAND2X1 NAND2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_8512_), .B(_8544_), .Y(_8545_) );
NAND2X1 NAND2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(module_1_H_18_), .Y(_8546_) );
AOI21X1 AOI21X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_8545_), .B(_8546_), .C(_8543_), .Y(_8547_) );
NAND2X1 NAND2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_19_), .B(_8517_), .Y(_8469_) );
NAND2X1 NAND2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_18_), .B(_8512_), .Y(_8470_) );
OAI21X1 OAI21X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_8543_), .B(_8470_), .C(_8469_), .Y(_8471_) );
AOI21X1 AOI21X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_8542_), .B(_8547_), .C(_8471_), .Y(_8472_) );
INVX1 INVX1_1178 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_23_), .Y(_8473_) );
INVX1 INVX1_1179 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_22_), .Y(_8474_) );
OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_8473_), .B(target[7]), .C(target[6]), .D(_8474_), .Y(_8475_) );
OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_8525_), .B(module_1_H_23_), .C(_8526_), .D(module_1_H_22_), .Y(_8476_) );
NOR2X1 NOR2X1_669 ( .gnd(gnd), .vdd(vdd), .A(_8475_), .B(_8476_), .Y(_8477_) );
NAND2X1 NAND2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_21_), .B(_8532_), .Y(_8478_) );
NAND2X1 NAND2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_20_), .B(_8533_), .Y(_8479_) );
AND2X2 AND2X2_186 ( .gnd(gnd), .vdd(vdd), .A(_8478_), .B(_8479_), .Y(_8480_) );
INVX1 INVX1_1180 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_20_), .Y(_8481_) );
NOR2X1 NOR2X1_670 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_21_), .B(_8532_), .Y(_8482_) );
AOI21X1 AOI21X1_1222 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_8481_), .C(_8482_), .Y(_8483_) );
NAND3X1 NAND3X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_8480_), .B(_8483_), .C(_8477_), .Y(_8484_) );
AOI21X1 AOI21X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_8478_), .B(_8479_), .C(_8482_), .Y(_8485_) );
AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_8525_), .B(module_1_H_23_), .C(_8526_), .D(module_1_H_22_), .Y(_8486_) );
NOR2X1 NOR2X1_671 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_23_), .B(_8525_), .Y(_8487_) );
AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_8525_), .B(module_1_H_15_), .C(_8526_), .D(module_1_H_14_), .Y(_8488_) );
NOR2X1 NOR2X1_672 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_15_), .B(_8525_), .Y(_8489_) );
OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_8486_), .B(_8487_), .C(_8488_), .D(_8489_), .Y(_8490_) );
AOI21X1 AOI21X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_8477_), .B(_8485_), .C(_8490_), .Y(_8491_) );
OAI21X1 OAI21X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_8472_), .B(_8484_), .C(_8491_), .Y(_8492_) );
NOR2X1 NOR2X1_673 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf3), .B(_8492__bF_buf1), .Y(module_1_comparador_target_hash_0_terminado) );
INVX1 INVX1_1181 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_0_), .Y(_8493_) );
NOR3X1 NOR3X1_243 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf2), .B(_8493_), .C(_8492__bF_buf3), .Y(bounty_24_) );
INVX1 INVX1_1182 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_1_), .Y(_8494_) );
NOR3X1 NOR3X1_244 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf4), .B(_8494_), .C(_8492__bF_buf4), .Y(bounty_25_) );
INVX1 INVX1_1183 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_2_), .Y(_8495_) );
NOR3X1 NOR3X1_245 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf3), .B(_8495_), .C(_8492__bF_buf1), .Y(bounty_26_) );
INVX1 INVX1_1184 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_3_), .Y(_8496_) );
NOR3X1 NOR3X1_246 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf4), .B(_8496_), .C(_8492__bF_buf4), .Y(bounty_27_) );
INVX1 INVX1_1185 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_4_), .Y(_8497_) );
NOR3X1 NOR3X1_247 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf0), .B(_8497_), .C(_8492__bF_buf0), .Y(bounty_28_) );
INVX1 INVX1_1186 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_5_), .Y(_8498_) );
NOR3X1 NOR3X1_248 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf4), .B(_8498_), .C(_8492__bF_buf4), .Y(bounty_29_) );
INVX1 INVX1_1187 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_6_), .Y(_8499_) );
NOR3X1 NOR3X1_249 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf4), .B(_8499_), .C(_8492__bF_buf4), .Y(bounty_30_) );
INVX1 INVX1_1188 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_7_), .Y(_8500_) );
NOR3X1 NOR3X1_250 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf0), .B(_8500_), .C(_8492__bF_buf0), .Y(bounty_31_) );
INVX1 INVX1_1189 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_8501_) );
NOR3X1 NOR3X1_251 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf1), .B(_8501_), .C(_8492__bF_buf2), .Y(bounty_32_) );
NOR3X1 NOR3X1_252 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf1), .B(_8506_), .C(_8492__bF_buf2), .Y(bounty_33_) );
NOR3X1 NOR3X1_253 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf1), .B(_8513_), .C(_8492__bF_buf2), .Y(bounty_34_) );
INVX1 INVX1_1190 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_8502_) );
NOR3X1 NOR3X1_254 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf1), .B(_8502_), .C(_8492__bF_buf2), .Y(bounty_35_) );
NOR3X1 NOR3X1_255 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf2), .B(_8530_), .C(_8492__bF_buf3), .Y(bounty_36_) );
NOR3X1 NOR3X1_256 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf4), .B(_8529_), .C(_8492__bF_buf4), .Y(bounty_37_) );
NOR3X1 NOR3X1_257 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf2), .B(_8523_), .C(_8492__bF_buf3), .Y(bounty_38_) );
NOR3X1 NOR3X1_258 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf2), .B(_8522_), .C(_8492__bF_buf3), .Y(bounty_39_) );
INVX1 INVX1_1191 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_16_), .Y(_8503_) );
NOR3X1 NOR3X1_259 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf3), .B(_8503_), .C(_8492__bF_buf1), .Y(bounty_40_) );
NOR3X1 NOR3X1_260 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf3), .B(_8540_), .C(_8492__bF_buf1), .Y(bounty_41_) );
NOR3X1 NOR3X1_261 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf3), .B(_8544_), .C(_8492__bF_buf1), .Y(bounty_42_) );
INVX1 INVX1_1192 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_19_), .Y(_8504_) );
NOR3X1 NOR3X1_262 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf1), .B(_8504_), .C(_8492__bF_buf2), .Y(bounty_43_) );
NOR3X1 NOR3X1_263 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf2), .B(_8481_), .C(_8492__bF_buf3), .Y(bounty_44_) );
INVX1 INVX1_1193 ( .gnd(gnd), .vdd(vdd), .A(module_1_H_21_), .Y(_8505_) );
NOR3X1 NOR3X1_264 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf0), .B(_8505_), .C(_8492__bF_buf0), .Y(bounty_45_) );
NOR3X1 NOR3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf0), .B(_8474_), .C(_8492__bF_buf0), .Y(bounty_46_) );
NOR3X1 NOR3X1_266 ( .gnd(gnd), .vdd(vdd), .A(_8539__bF_buf0), .B(_8473_), .C(_8492__bF_buf0), .Y(bounty_47_) );
INVX1 INVX1_1194 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf0_), .Y(_8548_) );
AOI21X1 AOI21X1_1225 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_24_), .B(_8548_), .C(bloque_datos_80_bF_buf0_), .Y(_8549_) );
OAI21X1 OAI21X1_1366 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_24_), .B(_8548_), .C(_8549_), .Y(module_1_W_136_) );
INVX1 INVX1_1195 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf1_), .Y(_8550_) );
AOI21X1 AOI21X1_1226 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_25_), .B(_8550_), .C(bloque_datos_81_bF_buf1_), .Y(_8551_) );
OAI21X1 OAI21X1_1367 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_25_), .B(_8550_), .C(_8551_), .Y(module_1_W_137_) );
INVX1 INVX1_1196 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf0_), .Y(_8552_) );
AOI21X1 AOI21X1_1227 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_26_), .B(_8552_), .C(bloque_datos_82_bF_buf0_), .Y(_8553_) );
OAI21X1 OAI21X1_1368 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_26_), .B(_8552_), .C(_8553_), .Y(module_1_W_138_) );
INVX1 INVX1_1197 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf0_), .Y(_8554_) );
AOI21X1 AOI21X1_1228 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_27_), .B(_8554_), .C(bloque_datos_83_bF_buf0_), .Y(_8555_) );
OAI21X1 OAI21X1_1369 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_27_), .B(_8554_), .C(_8555_), .Y(module_1_W_139_) );
INVX1 INVX1_1198 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf3_), .Y(_8556_) );
AOI21X1 AOI21X1_1229 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_28_), .B(_8556_), .C(bloque_datos_84_bF_buf0_), .Y(_8557_) );
OAI21X1 OAI21X1_1370 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_28_), .B(_8556_), .C(_8557_), .Y(module_1_W_140_) );
INVX1 INVX1_1199 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf3_), .Y(_8558_) );
AOI21X1 AOI21X1_1230 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_29_), .B(_8558_), .C(bloque_datos_85_bF_buf4_), .Y(_8559_) );
OAI21X1 OAI21X1_1371 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_29_), .B(_8558_), .C(_8559_), .Y(module_1_W_141_) );
INVX1 INVX1_1200 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf3_), .Y(_8560_) );
AOI21X1 AOI21X1_1231 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_30_), .B(_8560_), .C(bloque_datos_86_bF_buf0_), .Y(_8561_) );
OAI21X1 OAI21X1_1372 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_30_), .B(_8560_), .C(_8561_), .Y(module_1_W_142_) );
INVX1 INVX1_1201 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .Y(_8562_) );
AOI21X1 AOI21X1_1232 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_31_), .B(_8562_), .C(bloque_datos_87_bF_buf0_), .Y(_8563_) );
OAI21X1 OAI21X1_1373 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_31_), .B(_8562_), .C(_8563_), .Y(module_1_W_143_) );
INVX1 INVX1_1202 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf1_), .Y(_8564_) );
OR2X2 OR2X2_196 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_16_), .B(bloque_datos_24_bF_buf0_), .Y(_8565_) );
NAND2X1 NAND2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_16_), .B(bloque_datos_24_bF_buf4_), .Y(_8566_) );
NAND2X1 NAND2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_8566_), .B(_8565_), .Y(_8567_) );
NAND2X1 NAND2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_8564_), .B(_8567_), .Y(module_1_W_128_) );
INVX1 INVX1_1203 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf0_), .Y(_8568_) );
AOI21X1 AOI21X1_1233 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_17_), .B(_8568_), .C(bloque_datos_73_bF_buf2_), .Y(_8569_) );
OAI21X1 OAI21X1_1374 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_17_), .B(_8568_), .C(_8569_), .Y(module_1_W_129_) );
INVX1 INVX1_1204 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf1_), .Y(_8570_) );
OR2X2 OR2X2_197 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_18_), .B(bloque_datos_26_bF_buf2_), .Y(_8571_) );
NAND2X1 NAND2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_18_), .B(bloque_datos_26_bF_buf1_), .Y(_8572_) );
NAND2X1 NAND2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_8572_), .B(_8571_), .Y(_8573_) );
NAND2X1 NAND2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_8570_), .B(_8573_), .Y(module_1_W_130_) );
INVX1 INVX1_1205 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf4_), .Y(_8574_) );
OR2X2 OR2X2_198 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_19_), .B(bloque_datos_27_bF_buf4_), .Y(_8575_) );
NAND2X1 NAND2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_19_), .B(bloque_datos_27_bF_buf3_), .Y(_8576_) );
NAND2X1 NAND2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_8576_), .B(_8575_), .Y(_8577_) );
NAND2X1 NAND2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_8574_), .B(_8577_), .Y(module_1_W_131_) );
INVX2 INVX2_296 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf4_), .Y(_8578_) );
AOI21X1 AOI21X1_1234 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_20_), .B(_8578_), .C(bloque_datos_76_bF_buf0_), .Y(_8579_) );
OAI21X1 OAI21X1_1375 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_20_), .B(_8578_), .C(_8579_), .Y(module_1_W_132_) );
INVX2 INVX2_297 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf4_), .Y(_8580_) );
AOI21X1 AOI21X1_1235 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_21_), .B(_8580_), .C(bloque_datos_77_bF_buf0_), .Y(_8581_) );
OAI21X1 OAI21X1_1376 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_21_), .B(_8580_), .C(_8581_), .Y(module_1_W_133_) );
INVX2 INVX2_298 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf3_), .Y(_8582_) );
AOI21X1 AOI21X1_1236 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_22_), .B(_8582_), .C(bloque_datos_78_bF_buf0_), .Y(_8583_) );
OAI21X1 OAI21X1_1377 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_22_), .B(_8582_), .C(_8583_), .Y(module_1_W_134_) );
INVX1 INVX1_1206 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf1_), .Y(_8584_) );
AOI21X1 AOI21X1_1237 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_23_), .B(_8584_), .C(bloque_datos_79_bF_buf2_), .Y(_8585_) );
OAI21X1 OAI21X1_1378 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_23_), .B(_8584_), .C(_8585_), .Y(module_1_W_135_) );
INVX1 INVX1_1207 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(_8586_) );
INVX1 INVX1_1208 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf4_), .Y(_8587_) );
OAI21X1 OAI21X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_8586_), .B(bloque_datos_40_bF_buf0_), .C(_8587_), .Y(_8588_) );
AOI21X1 AOI21X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_8586_), .B(bloque_datos_40_bF_buf4_), .C(_8588_), .Y(_8589_) );
INVX1 INVX1_1209 ( .gnd(gnd), .vdd(vdd), .A(_8589_), .Y(module_1_W_144_) );
INVX1 INVX1_1210 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(_8590_) );
INVX1 INVX1_1211 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf1_), .Y(_8591_) );
OAI21X1 OAI21X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_8590_), .B(bloque_datos_41_bF_buf0_), .C(_8591_), .Y(_8592_) );
AOI21X1 AOI21X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_8590_), .B(bloque_datos_41_bF_buf3_), .C(_8592_), .Y(_8593_) );
INVX1 INVX1_1212 ( .gnd(gnd), .vdd(vdd), .A(_8593_), .Y(module_1_W_145_) );
INVX1 INVX1_1213 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf0_), .Y(_8594_) );
INVX1 INVX1_1214 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf4_), .Y(_8595_) );
OAI21X1 OAI21X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_8594_), .B(bloque_datos_42_bF_buf0_), .C(_8595_), .Y(_8596_) );
AOI21X1 AOI21X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_8594_), .B(bloque_datos_42_bF_buf3_), .C(_8596_), .Y(_8597_) );
INVX1 INVX1_1215 ( .gnd(gnd), .vdd(vdd), .A(_8597_), .Y(module_1_W_146_) );
INVX1 INVX1_1216 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf0_), .Y(_8598_) );
INVX1 INVX1_1217 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf3_), .Y(_8599_) );
OAI21X1 OAI21X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_8598_), .B(bloque_datos_43_bF_buf0_), .C(_8599_), .Y(_8600_) );
AOI21X1 AOI21X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_8598_), .B(bloque_datos_43_bF_buf3_), .C(_8600_), .Y(_8601_) );
INVX1 INVX1_1218 ( .gnd(gnd), .vdd(vdd), .A(_8601_), .Y(module_1_W_147_) );
INVX1 INVX1_1219 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf0_), .Y(_8602_) );
INVX1 INVX1_1220 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf0_), .Y(_8603_) );
OAI21X1 OAI21X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_8602_), .B(bloque_datos_44_bF_buf0_), .C(_8603_), .Y(_8604_) );
AOI21X1 AOI21X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_8602_), .B(bloque_datos_44_bF_buf4_), .C(_8604_), .Y(_8605_) );
INVX1 INVX1_1221 ( .gnd(gnd), .vdd(vdd), .A(_8605_), .Y(module_1_W_148_) );
INVX1 INVX1_1222 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf0_), .Y(_8606_) );
INVX1 INVX1_1223 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf0_), .Y(_8607_) );
OAI21X1 OAI21X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_8606_), .B(bloque_datos_45_bF_buf0_), .C(_8607_), .Y(_8608_) );
AOI21X1 AOI21X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_8606_), .B(bloque_datos_45_bF_buf4_), .C(_8608_), .Y(_8609_) );
INVX1 INVX1_1224 ( .gnd(gnd), .vdd(vdd), .A(_8609_), .Y(module_1_W_149_) );
INVX1 INVX1_1225 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf0_), .Y(_8610_) );
INVX1 INVX1_1226 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf0_), .Y(_8611_) );
OAI21X1 OAI21X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_8610_), .B(bloque_datos_46_bF_buf0_), .C(_8611_), .Y(_8612_) );
AOI21X1 AOI21X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_8610_), .B(bloque_datos_46_bF_buf4_), .C(_8612_), .Y(_8613_) );
INVX2 INVX2_299 ( .gnd(gnd), .vdd(vdd), .A(_8613_), .Y(module_1_W_150_) );
INVX1 INVX1_1227 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[7]), .Y(_8614_) );
INVX1 INVX1_1228 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf1_), .Y(_8615_) );
OAI21X1 OAI21X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_8614_), .B(bloque_datos_47_bF_buf2_), .C(_8615_), .Y(_8616_) );
AOI21X1 AOI21X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_8614_), .B(bloque_datos_47_bF_buf1_), .C(_8616_), .Y(_8617_) );
INVX2 INVX2_300 ( .gnd(gnd), .vdd(vdd), .A(_8617_), .Y(module_1_W_151_) );
AOI21X1 AOI21X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_8566_), .B(_8565_), .C(bloque_datos_72_bF_buf0_), .Y(_8618_) );
XNOR2X1 XNOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .B(bloque_datos_48_bF_buf0_), .Y(_8619_) );
NAND2X1 NAND2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_8619_), .B(_8618_), .Y(module_1_W_152_) );
XOR2X1 XOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .B(bloque_datos_49_bF_buf2_), .Y(_8620_) );
NOR2X1 NOR2X1_674 ( .gnd(gnd), .vdd(vdd), .A(_8620_), .B(module_1_W_129_), .Y(_8621_) );
INVX1 INVX1_1229 ( .gnd(gnd), .vdd(vdd), .A(_8621_), .Y(module_1_W_153_) );
AOI21X1 AOI21X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_8572_), .B(_8571_), .C(bloque_datos_74_bF_buf0_), .Y(_8622_) );
XNOR2X1 XNOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .B(bloque_datos_50_bF_buf0_), .Y(_8623_) );
NAND2X1 NAND2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_8623_), .B(_8622_), .Y(module_1_W_154_) );
AOI21X1 AOI21X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_8576_), .B(_8575_), .C(bloque_datos_75_bF_buf3_), .Y(_8624_) );
XNOR2X1 XNOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .B(bloque_datos_51_bF_buf4_), .Y(_8625_) );
NAND2X1 NAND2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_8625_), .B(_8624_), .Y(module_1_W_155_) );
INVX1 INVX1_1230 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_20_), .Y(_8626_) );
INVX1 INVX1_1231 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf4_), .Y(_8627_) );
OAI21X1 OAI21X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_8626_), .B(bloque_datos_28_bF_buf3_), .C(_8627_), .Y(_8628_) );
AOI21X1 AOI21X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_8626_), .B(bloque_datos_28_bF_buf2_), .C(_8628_), .Y(_8629_) );
AND2X2 AND2X2_187 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf3_), .B(bloque_datos_52_bF_buf0_), .Y(_8630_) );
NOR2X1 NOR2X1_675 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf2_), .B(bloque_datos_52_bF_buf4_), .Y(_8631_) );
OAI21X1 OAI21X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_8630_), .B(_8631_), .C(_8629_), .Y(module_1_W_156_) );
XOR2X1 XOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf0_), .B(bloque_datos_53_bF_buf3_), .Y(_8632_) );
NOR2X1 NOR2X1_676 ( .gnd(gnd), .vdd(vdd), .A(_8632_), .B(module_1_W_133_), .Y(_8633_) );
INVX1 INVX1_1232 ( .gnd(gnd), .vdd(vdd), .A(_8633_), .Y(module_1_W_157_) );
XOR2X1 XOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf0_), .B(bloque_datos_54_bF_buf3_), .Y(_8634_) );
NOR2X1 NOR2X1_677 ( .gnd(gnd), .vdd(vdd), .A(_8634_), .B(module_1_W_134_), .Y(_8635_) );
INVX1 INVX1_1233 ( .gnd(gnd), .vdd(vdd), .A(_8635_), .Y(module_1_W_158_) );
XOR2X1 XOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[15]), .B(bloque_datos[55]), .Y(_8636_) );
NOR2X1 NOR2X1_678 ( .gnd(gnd), .vdd(vdd), .A(_8636_), .B(module_1_W_135_), .Y(_8637_) );
INVX1 INVX1_1234 ( .gnd(gnd), .vdd(vdd), .A(_8637_), .Y(module_1_W_159_) );
XOR2X1 XOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_24_), .B(bloque_datos_32_bF_buf4_), .Y(_8638_) );
NOR2X1 NOR2X1_679 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf5_), .B(_8638_), .Y(_8639_) );
XNOR2X1 XNOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf0_), .B(bloque_datos_56_bF_buf0_), .Y(_8640_) );
NAND2X1 NAND2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_8640_), .B(_8639_), .Y(module_1_W_160_) );
INVX1 INVX1_1235 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_25_), .Y(_8641_) );
INVX1 INVX1_1236 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf0_), .Y(_8642_) );
OAI21X1 OAI21X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_8641_), .B(bloque_datos_33_bF_buf0_), .C(_8642_), .Y(_8643_) );
AOI21X1 AOI21X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_8641_), .B(bloque_datos_33_bF_buf3_), .C(_8643_), .Y(_8644_) );
XNOR2X1 XNOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .B(bloque_datos_57_bF_buf0_), .Y(_8645_) );
NAND2X1 NAND2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_8645_), .B(_8644_), .Y(module_1_W_161_) );
XOR2X1 XOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_26_), .B(bloque_datos_34_bF_buf4_), .Y(_8646_) );
NOR2X1 NOR2X1_680 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf4_), .B(_8646_), .Y(_8647_) );
XNOR2X1 XNOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .B(bloque_datos_58_bF_buf0_), .Y(_8648_) );
NAND2X1 NAND2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_8648_), .B(_8647_), .Y(module_1_W_162_) );
XOR2X1 XOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_27_), .B(bloque_datos_35_bF_buf4_), .Y(_8649_) );
NOR2X1 NOR2X1_681 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf5_), .B(_8649_), .Y(_8650_) );
XNOR2X1 XNOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf0_), .B(bloque_datos_59_bF_buf0_), .Y(_8651_) );
NAND2X1 NAND2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_8651_), .B(_8650_), .Y(module_1_W_163_) );
XOR2X1 XOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf0_), .B(bloque_datos_60_bF_buf3_), .Y(_8652_) );
NOR2X1 NOR2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_8652_), .B(module_1_W_140_), .Y(_8653_) );
INVX1 INVX1_1237 ( .gnd(gnd), .vdd(vdd), .A(_8653_), .Y(module_1_W_164_) );
XOR2X1 XOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf0_), .B(bloque_datos_61_bF_buf0_), .Y(_8654_) );
NOR2X1 NOR2X1_683 ( .gnd(gnd), .vdd(vdd), .A(_8654_), .B(module_1_W_141_), .Y(_8655_) );
INVX1 INVX1_1238 ( .gnd(gnd), .vdd(vdd), .A(_8655_), .Y(module_1_W_165_) );
XOR2X1 XOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf0_), .B(bloque_datos_62_bF_buf3_), .Y(_8656_) );
NOR2X1 NOR2X1_684 ( .gnd(gnd), .vdd(vdd), .A(_8656_), .B(module_1_W_142_), .Y(_8657_) );
INVX2 INVX2_301 ( .gnd(gnd), .vdd(vdd), .A(_8657_), .Y(module_1_W_166_) );
XOR2X1 XOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf0_), .B(bloque_datos[63]), .Y(_8658_) );
NOR2X1 NOR2X1_685 ( .gnd(gnd), .vdd(vdd), .A(_8658_), .B(module_1_W_143_), .Y(_8659_) );
INVX1 INVX1_1239 ( .gnd(gnd), .vdd(vdd), .A(_8659_), .Y(module_1_W_167_) );
XNOR2X1 XNOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf3_), .B(bloque_datos_64_bF_buf0_), .Y(_8660_) );
AND2X2 AND2X2_188 ( .gnd(gnd), .vdd(vdd), .A(_8589_), .B(_8660_), .Y(_8661_) );
INVX2 INVX2_302 ( .gnd(gnd), .vdd(vdd), .A(_8661_), .Y(module_1_W_168_) );
XNOR2X1 XNOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf3_), .B(bloque_datos_65_bF_buf0_), .Y(_8662_) );
AND2X2 AND2X2_189 ( .gnd(gnd), .vdd(vdd), .A(_8593_), .B(_8662_), .Y(_8663_) );
INVX1 INVX1_1240 ( .gnd(gnd), .vdd(vdd), .A(_8663_), .Y(module_1_W_169_) );
XNOR2X1 XNOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf0_), .B(bloque_datos_66_bF_buf0_), .Y(_8664_) );
AND2X2 AND2X2_190 ( .gnd(gnd), .vdd(vdd), .A(_8597_), .B(_8664_), .Y(_8665_) );
INVX1 INVX1_1241 ( .gnd(gnd), .vdd(vdd), .A(_8665_), .Y(module_1_W_170_) );
AND2X2 AND2X2_191 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf2_), .B(bloque_datos_67_bF_buf4_), .Y(_8666_) );
NOR2X1 NOR2X1_686 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf1_), .B(bloque_datos_67_bF_buf3_), .Y(_8667_) );
OAI21X1 OAI21X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_8666_), .B(_8667_), .C(_8601_), .Y(module_1_W_171_) );
INVX2 INVX2_303 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf3_), .Y(_8668_) );
NOR2X1 NOR2X1_687 ( .gnd(gnd), .vdd(vdd), .A(_8578_), .B(_8668_), .Y(_8669_) );
NOR2X1 NOR2X1_688 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf1_), .B(bloque_datos_68_bF_buf2_), .Y(_8670_) );
OAI21X1 OAI21X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_8669_), .B(_8670_), .C(_8605_), .Y(module_1_W_172_) );
INVX2 INVX2_304 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf3_), .Y(_8671_) );
NOR2X1 NOR2X1_689 ( .gnd(gnd), .vdd(vdd), .A(_8580_), .B(_8671_), .Y(_8672_) );
NOR2X1 NOR2X1_690 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf3_), .B(bloque_datos_69_bF_buf2_), .Y(_8673_) );
OAI21X1 OAI21X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_8672_), .B(_8673_), .C(_8609_), .Y(module_1_W_173_) );
INVX2 INVX2_305 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf3_), .Y(_8674_) );
NOR2X1 NOR2X1_691 ( .gnd(gnd), .vdd(vdd), .A(_8582_), .B(_8674_), .Y(_8675_) );
NOR2X1 NOR2X1_692 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf2_), .B(bloque_datos_70_bF_buf2_), .Y(_8676_) );
OAI21X1 OAI21X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_8675_), .B(_8676_), .C(_8613_), .Y(module_1_W_174_) );
XNOR2X1 XNOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf0_), .B(bloque_datos_71_bF_buf1_), .Y(_8677_) );
AND2X2 AND2X2_192 ( .gnd(gnd), .vdd(vdd), .A(_8617_), .B(_8677_), .Y(_8678_) );
INVX1 INVX1_1242 ( .gnd(gnd), .vdd(vdd), .A(_8678_), .Y(module_1_W_175_) );
XNOR2X1 XNOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf3_), .B(bloque_datos_72_bF_buf4_), .Y(_8679_) );
NAND3X1 NAND3X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_8619_), .B(_8679_), .C(_8618_), .Y(module_1_W_176_) );
INVX1 INVX1_1243 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_17_), .Y(_8680_) );
NAND2X1 NAND2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf2_), .B(_8680_), .Y(_8681_) );
AND2X2 AND2X2_193 ( .gnd(gnd), .vdd(vdd), .A(_8569_), .B(_8681_), .Y(_8682_) );
INVX1 INVX1_1244 ( .gnd(gnd), .vdd(vdd), .A(_8620_), .Y(_8683_) );
XNOR2X1 XNOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf2_), .B(bloque_datos_73_bF_buf1_), .Y(_8684_) );
NAND3X1 NAND3X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_8683_), .B(_8684_), .C(_8682_), .Y(module_1_W_177_) );
XNOR2X1 XNOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf3_), .B(bloque_datos_74_bF_buf4_), .Y(_8685_) );
NAND3X1 NAND3X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_8623_), .B(_8685_), .C(_8622_), .Y(module_1_W_178_) );
XNOR2X1 XNOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf3_), .B(bloque_datos_75_bF_buf2_), .Y(_8686_) );
NAND3X1 NAND3X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_8625_), .B(_8686_), .C(_8624_), .Y(module_1_W_179_) );
XOR2X1 XOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf2_), .B(bloque_datos_76_bF_buf3_), .Y(_8687_) );
NOR2X1 NOR2X1_693 ( .gnd(gnd), .vdd(vdd), .A(_8687_), .B(module_1_W_156_), .Y(_8688_) );
INVX1 INVX1_1245 ( .gnd(gnd), .vdd(vdd), .A(_8688_), .Y(module_1_W_180_) );
INVX1 INVX1_1246 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_21_), .Y(_8689_) );
INVX1 INVX1_1247 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf4_), .Y(_8690_) );
OAI21X1 OAI21X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_8689_), .B(bloque_datos_29_bF_buf2_), .C(_8690_), .Y(_8691_) );
AOI21X1 AOI21X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_8689_), .B(bloque_datos_29_bF_buf1_), .C(_8691_), .Y(_8692_) );
INVX1 INVX1_1248 ( .gnd(gnd), .vdd(vdd), .A(_8632_), .Y(_8693_) );
XNOR2X1 XNOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf2_), .B(bloque_datos_77_bF_buf3_), .Y(_8694_) );
NAND3X1 NAND3X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_8693_), .B(_8694_), .C(_8692_), .Y(module_1_W_181_) );
XNOR2X1 XNOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf2_), .B(bloque_datos_78_bF_buf4_), .Y(_8695_) );
AND2X2 AND2X2_194 ( .gnd(gnd), .vdd(vdd), .A(_8635_), .B(_8695_), .Y(_8696_) );
INVX2 INVX2_306 ( .gnd(gnd), .vdd(vdd), .A(_8696_), .Y(module_1_W_182_) );
XNOR2X1 XNOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .B(bloque_datos_79_bF_buf1_), .Y(_8697_) );
AND2X2 AND2X2_195 ( .gnd(gnd), .vdd(vdd), .A(_8637_), .B(_8697_), .Y(_8698_) );
INVX2 INVX2_307 ( .gnd(gnd), .vdd(vdd), .A(_8698_), .Y(module_1_W_183_) );
XNOR2X1 XNOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf4_), .B(bloque_datos_40_bF_buf3_), .Y(_8699_) );
NAND3X1 NAND3X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_8640_), .B(_8699_), .C(_8639_), .Y(module_1_W_184_) );
XNOR2X1 XNOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf4_), .B(bloque_datos_41_bF_buf2_), .Y(_8700_) );
NAND3X1 NAND3X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_8645_), .B(_8700_), .C(_8644_), .Y(module_1_W_185_) );
XNOR2X1 XNOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf3_), .B(bloque_datos_42_bF_buf2_), .Y(_8701_) );
NAND3X1 NAND3X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_8648_), .B(_8701_), .C(_8647_), .Y(module_1_W_186_) );
XNOR2X1 XNOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf4_), .B(bloque_datos_43_bF_buf2_), .Y(_8702_) );
NAND3X1 NAND3X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_8651_), .B(_8702_), .C(_8650_), .Y(module_1_W_187_) );
XNOR2X1 XNOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf4_), .B(bloque_datos_44_bF_buf3_), .Y(_8703_) );
AND2X2 AND2X2_196 ( .gnd(gnd), .vdd(vdd), .A(_8653_), .B(_8703_), .Y(_8704_) );
INVX1 INVX1_1249 ( .gnd(gnd), .vdd(vdd), .A(_8704_), .Y(module_1_W_188_) );
XNOR2X1 XNOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf3_), .B(bloque_datos_45_bF_buf3_), .Y(_8705_) );
AND2X2 AND2X2_197 ( .gnd(gnd), .vdd(vdd), .A(_8655_), .B(_8705_), .Y(_8706_) );
INVX1 INVX1_1250 ( .gnd(gnd), .vdd(vdd), .A(_8706_), .Y(module_1_W_189_) );
XNOR2X1 XNOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf4_), .B(bloque_datos_46_bF_buf3_), .Y(_8707_) );
AND2X2 AND2X2_198 ( .gnd(gnd), .vdd(vdd), .A(_8657_), .B(_8707_), .Y(_8708_) );
INVX1 INVX1_1251 ( .gnd(gnd), .vdd(vdd), .A(_8708_), .Y(module_1_W_190_) );
XNOR2X1 XNOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf3_), .B(bloque_datos_47_bF_buf0_), .Y(_8709_) );
AND2X2 AND2X2_199 ( .gnd(gnd), .vdd(vdd), .A(_8659_), .B(_8709_), .Y(_8710_) );
INVX1 INVX1_1252 ( .gnd(gnd), .vdd(vdd), .A(_8710_), .Y(module_1_W_191_) );
AND2X2 AND2X2_200 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf3_), .B(bloque_datos_48_bF_buf4_), .Y(_8711_) );
NOR2X1 NOR2X1_694 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf2_), .B(bloque_datos_48_bF_buf3_), .Y(_8712_) );
OAI21X1 OAI21X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_8711_), .B(_8712_), .C(_8661_), .Y(module_1_W_192_) );
AND2X2 AND2X2_201 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf0_), .B(bloque_datos_49_bF_buf1_), .Y(_8713_) );
NOR2X1 NOR2X1_695 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf3_), .B(bloque_datos_49_bF_buf0_), .Y(_8714_) );
OAI21X1 OAI21X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_8713_), .B(_8714_), .C(_8663_), .Y(module_1_W_193_) );
AND2X2 AND2X2_202 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf3_), .B(bloque_datos_50_bF_buf3_), .Y(_8715_) );
NOR2X1 NOR2X1_696 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf2_), .B(bloque_datos_50_bF_buf2_), .Y(_8716_) );
OAI21X1 OAI21X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_8715_), .B(_8716_), .C(_8665_), .Y(module_1_W_194_) );
OR2X2 OR2X2_199 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_171_), .B(bloque_datos_51_bF_buf3_), .Y(module_1_W_195_) );
NOR2X1 NOR2X1_697 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf3_), .B(module_1_W_172_), .Y(_8717_) );
INVX1 INVX1_1253 ( .gnd(gnd), .vdd(vdd), .A(_8717_), .Y(module_1_W_196_) );
NOR2X1 NOR2X1_698 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf2_), .B(module_1_W_173_), .Y(_8718_) );
INVX1 INVX1_1254 ( .gnd(gnd), .vdd(vdd), .A(_8718_), .Y(module_1_W_197_) );
OR2X2 OR2X2_200 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_174_), .B(bloque_datos_54_bF_buf2_), .Y(module_1_W_198_) );
XNOR2X1 XNOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf0_), .B(bloque_datos[55]), .Y(_8719_) );
NAND2X1 NAND2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_8678_), .Y(module_1_W_199_) );
NAND2X1 NAND2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf4_), .B(module_1_W_128_), .Y(_8720_) );
INVX1 INVX1_1255 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf3_), .Y(_8721_) );
NAND2X1 NAND2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_8721_), .B(_8618_), .Y(_8722_) );
AOI21X1 AOI21X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_8722_), .B(_8720_), .C(module_1_W_176_), .Y(_8723_) );
INVX2 INVX2_308 ( .gnd(gnd), .vdd(vdd), .A(_8723_), .Y(module_1_W_200_) );
NAND2X1 NAND2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf3_), .B(module_1_W_129_), .Y(_8724_) );
OR2X2 OR2X2_201 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_129_), .B(bloque_datos_57_bF_buf2_), .Y(_8725_) );
AOI21X1 AOI21X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_8724_), .B(_8725_), .C(module_1_W_177_), .Y(_8726_) );
INVX1 INVX1_1256 ( .gnd(gnd), .vdd(vdd), .A(_8726_), .Y(module_1_W_201_) );
NAND2X1 NAND2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf4_), .B(module_1_W_130_), .Y(_8727_) );
INVX1 INVX1_1257 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf3_), .Y(_8728_) );
NAND2X1 NAND2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_8728_), .B(_8622_), .Y(_8729_) );
AOI21X1 AOI21X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_8729_), .B(_8727_), .C(module_1_W_178_), .Y(_8730_) );
INVX1 INVX1_1258 ( .gnd(gnd), .vdd(vdd), .A(_8730_), .Y(module_1_W_202_) );
NAND2X1 NAND2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf4_), .B(module_1_W_131_), .Y(_8731_) );
INVX1 INVX1_1259 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf3_), .Y(_8732_) );
NAND2X1 NAND2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_8732_), .B(_8624_), .Y(_8733_) );
AOI21X1 AOI21X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_8733_), .B(_8731_), .C(module_1_W_179_), .Y(_8734_) );
INVX1 INVX1_1260 ( .gnd(gnd), .vdd(vdd), .A(_8734_), .Y(module_1_W_203_) );
XNOR2X1 XNOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_132_), .B(bloque_datos_60_bF_buf2_), .Y(_8735_) );
NAND2X1 NAND2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8688_), .Y(module_1_W_204_) );
NAND2X1 NAND2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf4_), .B(module_1_W_133_), .Y(_8736_) );
OR2X2 OR2X2_202 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_133_), .B(bloque_datos_61_bF_buf3_), .Y(_8737_) );
AOI21X1 AOI21X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_8737_), .C(module_1_W_181_), .Y(_8738_) );
INVX1 INVX1_1261 ( .gnd(gnd), .vdd(vdd), .A(_8738_), .Y(module_1_W_205_) );
INVX2 INVX2_309 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf2_), .Y(_8739_) );
NAND2X1 NAND2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_8739_), .B(_8696_), .Y(module_1_W_206_) );
INVX2 INVX2_310 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[63]), .Y(_8740_) );
NAND2X1 NAND2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_8740_), .B(_8698_), .Y(module_1_W_207_) );
OAI21X1 OAI21X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_8638_), .B(bloque_datos_80_bF_buf3_), .C(bloque_datos_64_bF_buf4_), .Y(_8741_) );
OR2X2 OR2X2_203 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_136_), .B(bloque_datos_64_bF_buf3_), .Y(_8742_) );
AOI21X1 AOI21X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_8741_), .B(_8742_), .C(module_1_W_184_), .Y(_8743_) );
INVX1 INVX1_1262 ( .gnd(gnd), .vdd(vdd), .A(_8743_), .Y(module_1_W_208_) );
NAND2X1 NAND2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_65_bF_buf3_), .B(module_1_W_137_), .Y(_8744_) );
OR2X2 OR2X2_204 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_137_), .B(bloque_datos_65_bF_buf2_), .Y(_8745_) );
AOI21X1 AOI21X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_8744_), .B(_8745_), .C(module_1_W_185_), .Y(_8746_) );
INVX1 INVX1_1263 ( .gnd(gnd), .vdd(vdd), .A(_8746_), .Y(module_1_W_209_) );
OAI21X1 OAI21X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(bloque_datos_82_bF_buf2_), .C(bloque_datos_66_bF_buf4_), .Y(_8747_) );
OR2X2 OR2X2_205 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_138_), .B(bloque_datos_66_bF_buf3_), .Y(_8748_) );
AOI21X1 AOI21X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_8747_), .B(_8748_), .C(module_1_W_186_), .Y(_8749_) );
INVX1 INVX1_1264 ( .gnd(gnd), .vdd(vdd), .A(_8749_), .Y(module_1_W_210_) );
OAI21X1 OAI21X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_8649_), .B(bloque_datos_83_bF_buf3_), .C(bloque_datos_67_bF_buf2_), .Y(_8750_) );
OR2X2 OR2X2_206 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_139_), .B(bloque_datos_67_bF_buf1_), .Y(_8751_) );
AOI21X1 AOI21X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_8750_), .B(_8751_), .C(module_1_W_187_), .Y(_8752_) );
INVX1 INVX1_1265 ( .gnd(gnd), .vdd(vdd), .A(_8752_), .Y(module_1_W_211_) );
NAND2X1 NAND2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_8668_), .B(_8704_), .Y(module_1_W_212_) );
NAND2X1 NAND2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_8671_), .B(_8706_), .Y(module_1_W_213_) );
NAND2X1 NAND2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_8674_), .B(_8708_), .Y(module_1_W_214_) );
INVX1 INVX1_1266 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf0_), .Y(_8753_) );
NAND2X1 NAND2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_8753_), .B(_8710_), .Y(module_1_W_215_) );
OR2X2 OR2X2_207 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_192_), .B(bloque_datos_72_bF_buf3_), .Y(module_1_W_216_) );
OR2X2 OR2X2_208 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_193_), .B(bloque_datos_73_bF_buf0_), .Y(module_1_W_217_) );
OR2X2 OR2X2_209 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_194_), .B(bloque_datos_74_bF_buf3_), .Y(module_1_W_218_) );
OR2X2 OR2X2_210 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_195_), .B(bloque_datos_75_bF_buf1_), .Y(module_1_W_219_) );
NAND2X1 NAND2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_8627_), .B(_8717_), .Y(module_1_W_220_) );
NAND2X1 NAND2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_8690_), .B(_8718_), .Y(module_1_W_221_) );
OR2X2 OR2X2_211 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_198_), .B(bloque_datos_78_bF_buf3_), .Y(module_1_W_222_) );
OR2X2 OR2X2_212 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_199_), .B(bloque_datos_79_bF_buf0_), .Y(module_1_W_223_) );
XNOR2X1 XNOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_152_), .B(bloque_datos_80_bF_buf2_), .Y(_8754_) );
NAND2X1 NAND2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_8723_), .B(_8754_), .Y(module_1_W_224_) );
OAI21X1 OAI21X1_1401 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_129_), .B(_8620_), .C(bloque_datos_81_bF_buf3_), .Y(_8755_) );
NAND3X1 NAND3X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_8642_), .B(_8683_), .C(_8682_), .Y(_8756_) );
NAND2X1 NAND2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_8755_), .B(_8756_), .Y(_8757_) );
NAND2X1 NAND2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_8726_), .Y(module_1_W_225_) );
XNOR2X1 XNOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_154_), .B(bloque_datos_82_bF_buf1_), .Y(_8758_) );
NAND2X1 NAND2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_8730_), .B(_8758_), .Y(module_1_W_226_) );
XNOR2X1 XNOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_155_), .B(bloque_datos_83_bF_buf2_), .Y(_8759_) );
NAND2X1 NAND2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_8734_), .B(_8759_), .Y(module_1_W_227_) );
INVX1 INVX1_1267 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf3_), .Y(_8760_) );
NAND3X1 NAND3X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_8760_), .B(_8735_), .C(_8688_), .Y(module_1_W_228_) );
OAI21X1 OAI21X1_1402 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_133_), .B(_8632_), .C(bloque_datos_85_bF_buf2_), .Y(_8761_) );
INVX1 INVX1_1268 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf1_), .Y(_8762_) );
NAND3X1 NAND3X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_8762_), .B(_8693_), .C(_8692_), .Y(_8763_) );
NAND2X1 NAND2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8763_), .Y(_8764_) );
NAND2X1 NAND2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8738_), .Y(module_1_W_229_) );
INVX1 INVX1_1269 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf3_), .Y(_8765_) );
NAND3X1 NAND3X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_8765_), .B(_8739_), .C(_8696_), .Y(module_1_W_230_) );
INVX1 INVX1_1270 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf2_), .Y(_8766_) );
NAND3X1 NAND3X1_1958 ( .gnd(gnd), .vdd(vdd), .A(_8766_), .B(_8740_), .C(_8698_), .Y(module_1_W_231_) );
AOI21X1 AOI21X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_8640_), .B(_8639_), .C(_8587_), .Y(_8767_) );
NOR2X1 NOR2X1_699 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf1_), .B(module_1_W_160_), .Y(_8768_) );
OAI21X1 OAI21X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_8768_), .B(_8767_), .C(_8743_), .Y(module_1_W_232_) );
AOI21X1 AOI21X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_8645_), .B(_8644_), .C(_8591_), .Y(_8769_) );
NOR2X1 NOR2X1_700 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf2_), .B(module_1_W_161_), .Y(_8770_) );
OAI21X1 OAI21X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_8769_), .B(_8770_), .C(_8746_), .Y(module_1_W_233_) );
AOI21X1 AOI21X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_8648_), .B(_8647_), .C(_8595_), .Y(_8771_) );
NOR2X1 NOR2X1_701 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf1_), .B(module_1_W_162_), .Y(_8772_) );
OAI21X1 OAI21X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_8772_), .B(_8771_), .C(_8749_), .Y(module_1_W_234_) );
AOI21X1 AOI21X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_8651_), .B(_8650_), .C(_8599_), .Y(_8773_) );
NOR2X1 NOR2X1_702 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf2_), .B(module_1_W_163_), .Y(_8774_) );
OAI21X1 OAI21X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_8774_), .B(_8773_), .C(_8752_), .Y(module_1_W_235_) );
NAND3X1 NAND3X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_8603_), .B(_8668_), .C(_8704_), .Y(module_1_W_236_) );
NAND3X1 NAND3X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_8607_), .B(_8671_), .C(_8706_), .Y(module_1_W_237_) );
NAND3X1 NAND3X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_8611_), .B(_8674_), .C(_8708_), .Y(module_1_W_238_) );
NAND3X1 NAND3X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_8615_), .B(_8753_), .C(_8710_), .Y(module_1_W_239_) );
OR2X2 OR2X2_213 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_192_), .B(module_1_W_128_), .Y(module_1_W_240_) );
OR2X2 OR2X2_214 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_193_), .B(module_1_W_129_), .Y(module_1_W_241_) );
OR2X2 OR2X2_215 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_194_), .B(module_1_W_130_), .Y(module_1_W_242_) );
OR2X2 OR2X2_216 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_195_), .B(module_1_W_131_), .Y(module_1_W_243_) );
NAND2X1 NAND2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_8629_), .B(_8717_), .Y(module_1_W_244_) );
NAND2X1 NAND2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_8692_), .B(_8718_), .Y(module_1_W_245_) );
OR2X2 OR2X2_217 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_198_), .B(module_1_W_134_), .Y(module_1_W_246_) );
OR2X2 OR2X2_218 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_199_), .B(module_1_W_135_), .Y(module_1_W_247_) );
XNOR2X1 XNOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_176_), .B(module_1_W_136_), .Y(_8775_) );
NAND3X1 NAND3X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_8723_), .B(_8754_), .C(_8775_), .Y(module_1_W_248_) );
NAND3X1 NAND3X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_8644_), .B(_8757_), .C(_8726_), .Y(module_1_W_249_) );
XNOR2X1 XNOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_178_), .B(module_1_W_138_), .Y(_8776_) );
NAND3X1 NAND3X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_8730_), .B(_8758_), .C(_8776_), .Y(module_1_W_250_) );
XNOR2X1 XNOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_179_), .B(module_1_W_139_), .Y(_8777_) );
NAND3X1 NAND3X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_8734_), .B(_8759_), .C(_8777_), .Y(module_1_W_251_) );
INVX1 INVX1_1271 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_140_), .Y(_8778_) );
NAND3X1 NAND3X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_8778_), .B(_8735_), .C(_8688_), .Y(module_1_W_252_) );
INVX1 INVX1_1272 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_141_), .Y(_8779_) );
NAND3X1 NAND3X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_8764_), .C(_8738_), .Y(module_1_W_253_) );
INVX1 INVX1_1273 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_142_), .Y(_8780_) );
NAND3X1 NAND3X1_1969 ( .gnd(gnd), .vdd(vdd), .A(_8739_), .B(_8780_), .C(_8696_), .Y(module_1_W_254_) );
INVX1 INVX1_1274 ( .gnd(gnd), .vdd(vdd), .A(module_1_W_143_), .Y(_8781_) );
NAND3X1 NAND3X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_8740_), .B(_8781_), .C(_8698_), .Y(module_1_W_255_) );
NAND3X1 NAND3X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_9014_), .B(_9015_), .C(_9016_), .Y(_9017_) );
NAND2X1 NAND2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_200_), .B(_8999_), .Y(_9018_) );
OR2X2 OR2X2_219 ( .gnd(gnd), .vdd(vdd), .A(_8999_), .B(module_2_W_200_), .Y(_9019_) );
NAND2X1 NAND2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_9018_), .B(_9019_), .Y(_9020_) );
NAND3X1 NAND3X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_9017_), .B(_9020_), .C(_9012_), .Y(_9021_) );
NAND2X1 NAND2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_9017_), .B(_9012_), .Y(_9022_) );
INVX2 INVX2_311 ( .gnd(gnd), .vdd(vdd), .A(_9020_), .Y(_9023_) );
AOI21X1 AOI21X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_9022_), .C(_11005_), .Y(_9024_) );
NAND3X1 NAND3X1_1973 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_228_), .B(_9021_), .C(_9024_), .Y(_9025_) );
INVX1 INVX1_1275 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_228_), .Y(_9026_) );
AOI21X1 AOI21X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_9015_), .B(_9016_), .C(_9014_), .Y(_9027_) );
NAND3X1 NAND3X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_12434_), .B(_9007_), .C(_9004_), .Y(_9028_) );
NAND3X1 NAND3X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_12437_), .B(_9009_), .C(_9010_), .Y(_9029_) );
AOI21X1 AOI21X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_9028_), .B(_9029_), .C(_12490_), .Y(_9030_) );
OAI21X1 OAI21X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_9027_), .B(_9030_), .C(_9023_), .Y(_9031_) );
NAND3X1 NAND3X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_10994_), .B(_9021_), .C(_9031_), .Y(_9032_) );
NAND2X1 NAND2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_9026_), .B(_9032_), .Y(_9033_) );
AOI21X1 AOI21X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_9033_), .B(_9025_), .C(_12446_), .Y(_9034_) );
INVX1 INVX1_1276 ( .gnd(gnd), .vdd(vdd), .A(_12446_), .Y(_9035_) );
NAND2X1 NAND2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_228_), .B(_9032_), .Y(_9036_) );
NAND3X1 NAND3X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_9026_), .B(_9021_), .C(_9024_), .Y(_9037_) );
AOI21X1 AOI21X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_9036_), .B(_9037_), .C(_9035_), .Y(_9038_) );
OAI21X1 OAI21X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_9034_), .B(_9038_), .C(_12488_), .Y(_9039_) );
OAI21X1 OAI21X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_12452_), .B(_12454_), .C(_12447_), .Y(_9040_) );
NAND3X1 NAND3X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_9035_), .B(_9036_), .C(_9037_), .Y(_9041_) );
NAND3X1 NAND3X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_12446_), .B(_9033_), .C(_9025_), .Y(_9042_) );
NAND3X1 NAND3X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(_9041_), .C(_9042_), .Y(_9043_) );
NAND2X1 NAND2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_216_), .B(_9020_), .Y(_9044_) );
OR2X2 OR2X2_220 ( .gnd(gnd), .vdd(vdd), .A(_9020_), .B(module_2_W_216_), .Y(_9045_) );
NAND2X1 NAND2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_9044_), .B(_9045_), .Y(_9046_) );
NAND3X1 NAND3X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_9043_), .B(_9046_), .C(_9039_), .Y(_9047_) );
AOI21X1 AOI21X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_9041_), .B(_9042_), .C(_9040_), .Y(_9048_) );
NOR3X1 NOR3X1_267 ( .gnd(gnd), .vdd(vdd), .A(_9034_), .B(_9038_), .C(_12488_), .Y(_9049_) );
INVX2 INVX2_312 ( .gnd(gnd), .vdd(vdd), .A(_9046_), .Y(_9050_) );
OAI21X1 OAI21X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_9049_), .B(_9048_), .C(_9050_), .Y(_9051_) );
NAND3X1 NAND3X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_12239_), .B(_9047_), .C(_9051_), .Y(_9052_) );
NAND2X1 NAND2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_244_), .B(_9052_), .Y(_9053_) );
INVX1 INVX1_1277 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_244_), .Y(_9054_) );
NAND2X1 NAND2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_9043_), .B(_9039_), .Y(_9055_) );
AOI21X1 AOI21X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_9050_), .B(_9055_), .C(_12240_), .Y(_9056_) );
NAND3X1 NAND3X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_9054_), .B(_9047_), .C(_9056_), .Y(_9057_) );
NAND3X1 NAND3X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_12487_), .B(_9057_), .C(_9053_), .Y(_9058_) );
NAND3X1 NAND3X1_1985 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_244_), .B(_9047_), .C(_9056_), .Y(_9059_) );
NAND2X1 NAND2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_9054_), .B(_9052_), .Y(_9060_) );
NAND3X1 NAND3X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_12459_), .B(_9059_), .C(_9060_), .Y(_9061_) );
AOI21X1 AOI21X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_9058_), .B(_9061_), .C(_12486_), .Y(_9062_) );
NOR2X1 NOR2X1_703 ( .gnd(gnd), .vdd(vdd), .A(_12235_), .B(_12460_), .Y(_9063_) );
AOI21X1 AOI21X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_12250_), .B(_12463_), .C(_9063_), .Y(_9064_) );
AOI21X1 AOI21X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_9059_), .B(_9060_), .C(_12459_), .Y(_9065_) );
AOI21X1 AOI21X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_9057_), .B(_9053_), .C(_12487_), .Y(_9066_) );
NOR3X1 NOR3X1_268 ( .gnd(gnd), .vdd(vdd), .A(_9065_), .B(_9064_), .C(_9066_), .Y(_9067_) );
NOR2X1 NOR2X1_704 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_232_), .B(_9050_), .Y(_9068_) );
AND2X2 AND2X2_203 ( .gnd(gnd), .vdd(vdd), .A(_9050_), .B(module_2_W_232_), .Y(_9069_) );
NOR2X1 NOR2X1_705 ( .gnd(gnd), .vdd(vdd), .A(_9068_), .B(_9069_), .Y(_9070_) );
OAI21X1 OAI21X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_9067_), .B(_9062_), .C(_9070_), .Y(_9071_) );
OAI21X1 OAI21X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_9065_), .B(_9066_), .C(_9064_), .Y(_9072_) );
NAND3X1 NAND3X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_9058_), .B(_9061_), .C(_12486_), .Y(_9073_) );
INVX2 INVX2_313 ( .gnd(gnd), .vdd(vdd), .A(_9070_), .Y(_9074_) );
NAND3X1 NAND3X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_9074_), .B(_9073_), .C(_9072_), .Y(_9075_) );
NAND2X1 NAND2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_9075_), .B(_9071_), .Y(_9076_) );
XNOR2X1 XNOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_9076_), .B(_12483_), .Y(module_2_H_4_) );
NAND3X1 NAND3X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_12483_), .B(_9075_), .C(_9071_), .Y(_9077_) );
NOR2X1 NOR2X1_706 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_216_), .B(_9023_), .Y(_9078_) );
NOR2X1 NOR2X1_707 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_200_), .B(_9000_), .Y(_9079_) );
NOR2X1 NOR2X1_708 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_184_), .B(_8975_), .Y(_9080_) );
INVX1 INVX1_1278 ( .gnd(gnd), .vdd(vdd), .A(_8953_), .Y(_9081_) );
NOR2X1 NOR2X1_709 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_168_), .B(_9081_), .Y(_9082_) );
NOR2X1 NOR2X1_710 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_152_), .B(_8931_), .Y(_9083_) );
INVX1 INVX1_1279 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_153_), .Y(_9084_) );
NOR2X1 NOR2X1_711 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_136_), .B(_8908_), .Y(_9085_) );
INVX1 INVX1_1280 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_137_), .Y(_9086_) );
INVX1 INVX1_1281 ( .gnd(gnd), .vdd(vdd), .A(_8878_), .Y(_9087_) );
NOR2X1 NOR2X1_712 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf0_), .B(_9087_), .Y(_9088_) );
INVX1 INVX1_1282 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf1_), .Y(_9089_) );
INVX1 INVX1_1283 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_73_bF_buf3_), .Y(_9090_) );
NOR2X1 NOR2X1_713 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf2_), .B(_8828_), .Y(_9091_) );
NOR2X1 NOR2X1_714 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf2_), .B(_8803_), .Y(_9092_) );
NOR2X1 NOR2X1_715 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf2_), .B(_12589_), .Y(_9093_) );
NOR2X1 NOR2X1_716 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .B(_12564_), .Y(_9094_) );
INVX1 INVX1_1284 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_25_), .Y(_9095_) );
INVX2 INVX2_314 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_9_), .Y(_9096_) );
NOR2X1 NOR2X1_717 ( .gnd(gnd), .vdd(vdd), .A(_9095_), .B(_9096_), .Y(_9097_) );
NOR2X1 NOR2X1_718 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_25_), .B(module_2_W_9_), .Y(_9098_) );
NOR2X1 NOR2X1_719 ( .gnd(gnd), .vdd(vdd), .A(_9098_), .B(_9097_), .Y(_9099_) );
NOR2X1 NOR2X1_720 ( .gnd(gnd), .vdd(vdd), .A(_12562_), .B(_9099_), .Y(_9100_) );
AND2X2 AND2X2_204 ( .gnd(gnd), .vdd(vdd), .A(_9099_), .B(_12562_), .Y(_9101_) );
NOR2X1 NOR2X1_721 ( .gnd(gnd), .vdd(vdd), .A(_9100_), .B(_9101_), .Y(_9102_) );
NOR2X1 NOR2X1_722 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .B(_9102_), .Y(_9103_) );
INVX1 INVX1_1285 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .Y(_9104_) );
OR2X2 OR2X2_221 ( .gnd(gnd), .vdd(vdd), .A(_9101_), .B(_9100_), .Y(_9105_) );
NOR2X1 NOR2X1_723 ( .gnd(gnd), .vdd(vdd), .A(_9104_), .B(_9105_), .Y(_9106_) );
OAI21X1 OAI21X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_9106_), .B(_9103_), .C(_9094_), .Y(_9107_) );
OR2X2 OR2X2_222 ( .gnd(gnd), .vdd(vdd), .A(_9106_), .B(_9103_), .Y(_9108_) );
OR2X2 OR2X2_223 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_9094_), .Y(_9109_) );
AND2X2 AND2X2_205 ( .gnd(gnd), .vdd(vdd), .A(_9109_), .B(_9107_), .Y(_9110_) );
NOR2X1 NOR2X1_724 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf1_), .B(_9110_), .Y(_9111_) );
AND2X2 AND2X2_206 ( .gnd(gnd), .vdd(vdd), .A(_9110_), .B(bloque_datos_25_bF_buf0_), .Y(_9112_) );
OAI21X1 OAI21X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_9111_), .C(_9093_), .Y(_9113_) );
OR2X2 OR2X2_224 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_9111_), .Y(_9114_) );
OR2X2 OR2X2_225 ( .gnd(gnd), .vdd(vdd), .A(_9114_), .B(_9093_), .Y(_9115_) );
AND2X2 AND2X2_207 ( .gnd(gnd), .vdd(vdd), .A(_9115_), .B(_9113_), .Y(_9116_) );
NOR2X1 NOR2X1_725 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf1_), .B(_9116_), .Y(_9117_) );
INVX1 INVX1_1286 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf0_), .Y(_9118_) );
NAND2X1 NAND2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_9113_), .B(_9115_), .Y(_9119_) );
NOR2X1 NOR2X1_726 ( .gnd(gnd), .vdd(vdd), .A(_9118_), .B(_9119_), .Y(_9120_) );
OAI21X1 OAI21X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_9117_), .B(_9120_), .C(_9092_), .Y(_9121_) );
OR2X2 OR2X2_226 ( .gnd(gnd), .vdd(vdd), .A(_9117_), .B(_9120_), .Y(_9122_) );
OR2X2 OR2X2_227 ( .gnd(gnd), .vdd(vdd), .A(_9122_), .B(_9092_), .Y(_9123_) );
AND2X2 AND2X2_208 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_9121_), .Y(_9124_) );
NOR2X1 NOR2X1_727 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf1_), .B(_9124_), .Y(_9125_) );
INVX1 INVX1_1287 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf0_), .Y(_9126_) );
NAND2X1 NAND2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_9121_), .B(_9123_), .Y(_9127_) );
NOR2X1 NOR2X1_728 ( .gnd(gnd), .vdd(vdd), .A(_9126_), .B(_9127_), .Y(_9128_) );
OAI21X1 OAI21X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_9125_), .B(_9128_), .C(_9091_), .Y(_9129_) );
OR2X2 OR2X2_228 ( .gnd(gnd), .vdd(vdd), .A(_9125_), .B(_9128_), .Y(_9130_) );
OR2X2 OR2X2_229 ( .gnd(gnd), .vdd(vdd), .A(_9130_), .B(_9091_), .Y(_9131_) );
NAND2X1 NAND2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_9129_), .B(_9131_), .Y(_9132_) );
NAND2X1 NAND2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_9090_), .B(_9132_), .Y(_9133_) );
OR2X2 OR2X2_230 ( .gnd(gnd), .vdd(vdd), .A(_9132_), .B(_9090_), .Y(_9134_) );
NAND2X1 NAND2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_9133_), .B(_9134_), .Y(_9135_) );
NAND2X1 NAND2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_8875_), .B(_9135_), .Y(_9136_) );
OR2X2 OR2X2_231 ( .gnd(gnd), .vdd(vdd), .A(_9135_), .B(_8875_), .Y(_9137_) );
NAND2X1 NAND2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_9136_), .B(_9137_), .Y(_9138_) );
NAND2X1 NAND2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_9138_), .Y(_9139_) );
OR2X2 OR2X2_232 ( .gnd(gnd), .vdd(vdd), .A(_9138_), .B(_9089_), .Y(_9140_) );
NAND2X1 NAND2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_9139_), .B(_9140_), .Y(_9141_) );
NAND2X1 NAND2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_9088_), .B(_9141_), .Y(_9142_) );
NOR2X1 NOR2X1_729 ( .gnd(gnd), .vdd(vdd), .A(_9088_), .B(_9141_), .Y(_9143_) );
INVX1 INVX1_1288 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .Y(_9144_) );
NAND2X1 NAND2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_9142_), .B(_9144_), .Y(_9145_) );
NAND2X1 NAND2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_9086_), .B(_9145_), .Y(_9146_) );
INVX2 INVX2_315 ( .gnd(gnd), .vdd(vdd), .A(_9145_), .Y(_9147_) );
NAND2X1 NAND2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_137_), .B(_9147_), .Y(_9148_) );
NAND2X1 NAND2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_9146_), .B(_9148_), .Y(_9149_) );
NAND2X1 NAND2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_9085_), .B(_9149_), .Y(_9150_) );
NOR2X1 NOR2X1_730 ( .gnd(gnd), .vdd(vdd), .A(_9085_), .B(_9149_), .Y(_9151_) );
INVX1 INVX1_1289 ( .gnd(gnd), .vdd(vdd), .A(_9151_), .Y(_9152_) );
NAND2X1 NAND2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_9150_), .B(_9152_), .Y(_9153_) );
NAND2X1 NAND2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_9084_), .B(_9153_), .Y(_9154_) );
NOR2X1 NOR2X1_731 ( .gnd(gnd), .vdd(vdd), .A(_9084_), .B(_9153_), .Y(_9155_) );
INVX1 INVX1_1290 ( .gnd(gnd), .vdd(vdd), .A(_9155_), .Y(_9156_) );
NAND2X1 NAND2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_9154_), .B(_9156_), .Y(_9157_) );
NAND2X1 NAND2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_9083_), .B(_9157_), .Y(_9158_) );
NOR2X1 NOR2X1_732 ( .gnd(gnd), .vdd(vdd), .A(_9083_), .B(_9157_), .Y(_9159_) );
INVX1 INVX1_1291 ( .gnd(gnd), .vdd(vdd), .A(_9159_), .Y(_9160_) );
NAND2X1 NAND2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_9158_), .B(_9160_), .Y(_9161_) );
INVX2 INVX2_316 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .Y(_9162_) );
NOR2X1 NOR2X1_733 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_169_), .B(_9162_), .Y(_9163_) );
NAND2X1 NAND2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_169_), .B(_9162_), .Y(_9164_) );
INVX2 INVX2_317 ( .gnd(gnd), .vdd(vdd), .A(_9164_), .Y(_9165_) );
OAI21X1 OAI21X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_9165_), .B(_9163_), .C(_9082_), .Y(_9166_) );
NOR2X1 NOR2X1_734 ( .gnd(gnd), .vdd(vdd), .A(_9163_), .B(_9165_), .Y(_9167_) );
OAI21X1 OAI21X1_1418 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_168_), .B(_9081_), .C(_9167_), .Y(_9168_) );
NAND2X1 NAND2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_9166_), .B(_9168_), .Y(_9169_) );
INVX2 INVX2_318 ( .gnd(gnd), .vdd(vdd), .A(_9169_), .Y(_9170_) );
NOR2X1 NOR2X1_735 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_185_), .B(_9170_), .Y(_9171_) );
NAND2X1 NAND2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_185_), .B(_9170_), .Y(_9172_) );
INVX2 INVX2_319 ( .gnd(gnd), .vdd(vdd), .A(_9172_), .Y(_9173_) );
OAI21X1 OAI21X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_9173_), .B(_9171_), .C(_9080_), .Y(_9174_) );
NOR2X1 NOR2X1_736 ( .gnd(gnd), .vdd(vdd), .A(_9171_), .B(_9173_), .Y(_9175_) );
OAI21X1 OAI21X1_1420 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_184_), .B(_8975_), .C(_9175_), .Y(_9176_) );
NAND2X1 NAND2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_9174_), .B(_9176_), .Y(_9177_) );
INVX2 INVX2_320 ( .gnd(gnd), .vdd(vdd), .A(_9177_), .Y(_9178_) );
NOR2X1 NOR2X1_737 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_201_), .B(_9178_), .Y(_9179_) );
NAND2X1 NAND2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_201_), .B(_9178_), .Y(_9180_) );
INVX2 INVX2_321 ( .gnd(gnd), .vdd(vdd), .A(_9180_), .Y(_9181_) );
OAI21X1 OAI21X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_9181_), .B(_9179_), .C(_9079_), .Y(_9182_) );
NOR2X1 NOR2X1_738 ( .gnd(gnd), .vdd(vdd), .A(_9179_), .B(_9181_), .Y(_9183_) );
OAI21X1 OAI21X1_1422 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_200_), .B(_9000_), .C(_9183_), .Y(_9184_) );
NAND2X1 NAND2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_9182_), .B(_9184_), .Y(_9185_) );
INVX2 INVX2_322 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .Y(_9186_) );
NOR2X1 NOR2X1_739 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_217_), .B(_9186_), .Y(_9187_) );
NAND2X1 NAND2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_217_), .B(_9186_), .Y(_9188_) );
INVX2 INVX2_323 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .Y(_9189_) );
OAI21X1 OAI21X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_9189_), .B(_9187_), .C(_9078_), .Y(_9190_) );
NOR2X1 NOR2X1_740 ( .gnd(gnd), .vdd(vdd), .A(_9187_), .B(_9189_), .Y(_9191_) );
OAI21X1 OAI21X1_1424 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_216_), .B(_9023_), .C(_9191_), .Y(_9192_) );
NAND2X1 NAND2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_9190_), .B(_9192_), .Y(_9193_) );
INVX2 INVX2_324 ( .gnd(gnd), .vdd(vdd), .A(_9193_), .Y(_9194_) );
NOR2X1 NOR2X1_741 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_233_), .B(_9194_), .Y(_9195_) );
NAND2X1 NAND2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_233_), .B(_9194_), .Y(_9196_) );
INVX2 INVX2_325 ( .gnd(gnd), .vdd(vdd), .A(_9196_), .Y(_9197_) );
OAI21X1 OAI21X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_9195_), .C(_9068_), .Y(_9198_) );
NOR2X1 NOR2X1_742 ( .gnd(gnd), .vdd(vdd), .A(_9195_), .B(_9197_), .Y(_9199_) );
OAI21X1 OAI21X1_1426 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_232_), .B(_9050_), .C(_9199_), .Y(_9200_) );
NAND2X1 NAND2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_9198_), .B(_9200_), .Y(_9201_) );
OAI21X1 OAI21X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_9066_), .B(_9064_), .C(_9058_), .Y(_9202_) );
INVX1 INVX1_1292 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_245_), .Y(_9203_) );
AOI21X1 AOI21X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(_9042_), .C(_9034_), .Y(_9204_) );
INVX2 INVX2_326 ( .gnd(gnd), .vdd(vdd), .A(_9036_), .Y(_9205_) );
INVX1 INVX1_1293 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_229_), .Y(_9206_) );
AOI21X1 AOI21X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_9014_), .B(_9016_), .C(_9008_), .Y(_9207_) );
INVX2 INVX2_327 ( .gnd(gnd), .vdd(vdd), .A(_9009_), .Y(_9208_) );
INVX1 INVX1_1294 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_213_), .Y(_9209_) );
AOI21X1 AOI21X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_8994_), .B(_8992_), .C(_8984_), .Y(_9210_) );
INVX2 INVX2_328 ( .gnd(gnd), .vdd(vdd), .A(_8988_), .Y(_9211_) );
INVX1 INVX1_1295 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_197_), .Y(_9212_) );
AOI21X1 AOI21X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_8968_), .B(_8966_), .C(_8961_), .Y(_9213_) );
INVX2 INVX2_329 ( .gnd(gnd), .vdd(vdd), .A(_8962_), .Y(_9214_) );
INVX1 INVX1_1296 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_181_), .Y(_9215_) );
AOI21X1 AOI21X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_12496_), .B(_8949_), .C(_8942_), .Y(_9216_) );
INVX2 INVX2_330 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .Y(_9217_) );
INVX1 INVX1_1297 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_165_), .Y(_9218_) );
INVX1 INVX1_1298 ( .gnd(gnd), .vdd(vdd), .A(_9153_), .Y(_9219_) );
AOI21X1 AOI21X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_8922_), .B(_8924_), .C(_8917_), .Y(_9220_) );
INVX1 INVX1_1299 ( .gnd(gnd), .vdd(vdd), .A(_8918_), .Y(_9221_) );
INVX1 INVX1_1300 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_149_), .Y(_9222_) );
AOI21X1 AOI21X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_8894_), .B(_12499_), .C(_8904_), .Y(_9223_) );
AOI21X1 AOI21X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_8867_), .B(_8868_), .C(_12501_), .Y(_9224_) );
AOI21X1 AOI21X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8873_), .C(_9224_), .Y(_9225_) );
NOR3X1 NOR3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_8835_), .B(_12353_), .C(_8839_), .Y(_9226_) );
OAI21X1 OAI21X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_9226_), .B(_12503_), .C(_8848_), .Y(_9227_) );
AOI21X1 AOI21X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_8817_), .B(_8818_), .C(_12507_), .Y(_9228_) );
AOI21X1 AOI21X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_8823_), .B(_8821_), .C(_9228_), .Y(_9229_) );
AOI21X1 AOI21X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_8792_), .B(_8793_), .C(_12511_), .Y(_9230_) );
AOI21X1 AOI21X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_8798_), .B(_8796_), .C(_9230_), .Y(_9231_) );
INVX1 INVX1_1301 ( .gnd(gnd), .vdd(vdd), .A(_12582_), .Y(_9232_) );
AOI21X1 AOI21X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_12581_), .B(_12583_), .C(_9232_), .Y(_9233_) );
INVX1 INVX1_1302 ( .gnd(gnd), .vdd(vdd), .A(_12558_), .Y(_9234_) );
AOI21X1 AOI21X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_12559_), .B(_12557_), .C(_9234_), .Y(_9235_) );
AOI21X1 AOI21X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_12531_), .B(_12530_), .C(_12290_), .Y(_9236_) );
NOR2X1 NOR2X1_743 ( .gnd(gnd), .vdd(vdd), .A(_9236_), .B(_12542_), .Y(_9237_) );
INVX1 INVX1_1303 ( .gnd(gnd), .vdd(vdd), .A(_12530_), .Y(_9238_) );
NOR2X1 NOR2X1_744 ( .gnd(gnd), .vdd(vdd), .A(_11389_), .B(_11378_), .Y(_9239_) );
INVX2 INVX2_331 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_5_), .Y(_9240_) );
XNOR2X1 XNOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_12522_), .B(_9240_), .Y(_9241_) );
NAND2X1 NAND2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_9239_), .B(_9241_), .Y(_9242_) );
INVX1 INVX1_1304 ( .gnd(gnd), .vdd(vdd), .A(_9239_), .Y(_9243_) );
NOR2X1 NOR2X1_745 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_5_), .B(_12522_), .Y(_9244_) );
NOR2X1 NOR2X1_746 ( .gnd(gnd), .vdd(vdd), .A(_9240_), .B(_12519_), .Y(_9245_) );
OAI21X1 OAI21X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_9245_), .B(_9244_), .C(_9243_), .Y(_9246_) );
NAND3X1 NAND3X1_1990 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_21_), .B(_9242_), .C(_9246_), .Y(_9247_) );
INVX1 INVX1_1305 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_21_), .Y(_9248_) );
OAI21X1 OAI21X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_9245_), .B(_9244_), .C(_9239_), .Y(_9249_) );
OAI21X1 OAI21X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_11378_), .B(_11389_), .C(_9241_), .Y(_9250_) );
NAND3X1 NAND3X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_9248_), .B(_9250_), .C(_9249_), .Y(_9251_) );
NAND3X1 NAND3X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_9238_), .B(_9247_), .C(_9251_), .Y(_9252_) );
NAND3X1 NAND3X1_1993 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_21_), .B(_9250_), .C(_9249_), .Y(_9253_) );
NAND3X1 NAND3X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_9248_), .B(_9242_), .C(_9246_), .Y(_9254_) );
NAND3X1 NAND3X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_12530_), .B(_9254_), .C(_9253_), .Y(_9255_) );
AND2X2 AND2X2_209 ( .gnd(gnd), .vdd(vdd), .A(_9252_), .B(_9255_), .Y(_9256_) );
NAND2X1 NAND2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_9256_), .B(_9237_), .Y(_9257_) );
NAND2X1 NAND2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_9255_), .B(_9252_), .Y(_9258_) );
OAI21X1 OAI21X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_9236_), .B(_12542_), .C(_9258_), .Y(_9259_) );
XNOR2X1 XNOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_11465_), .B(module_2_W_9_), .Y(_9260_) );
NAND3X1 NAND3X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(_9259_), .C(_9257_), .Y(_9261_) );
NAND2X1 NAND2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_12529_), .B(_12533_), .Y(_9262_) );
NOR2X1 NOR2X1_747 ( .gnd(gnd), .vdd(vdd), .A(_9258_), .B(_9262_), .Y(_9263_) );
NOR2X1 NOR2X1_748 ( .gnd(gnd), .vdd(vdd), .A(_9256_), .B(_9237_), .Y(_9264_) );
INVX1 INVX1_1306 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .Y(_9265_) );
OAI21X1 OAI21X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_9264_), .B(_9263_), .C(_9265_), .Y(_9266_) );
NAND3X1 NAND3X1_1997 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf3_), .B(_9261_), .C(_9266_), .Y(_9267_) );
INVX1 INVX1_1307 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf2_), .Y(_9268_) );
NAND3X1 NAND3X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_9265_), .B(_9259_), .C(_9257_), .Y(_9269_) );
OAI21X1 OAI21X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_9264_), .B(_9263_), .C(_9260_), .Y(_9270_) );
NAND3X1 NAND3X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .B(_9269_), .C(_9270_), .Y(_9271_) );
NAND3X1 NAND3X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_12545_), .B(_9267_), .C(_9271_), .Y(_9272_) );
NAND3X1 NAND3X1_2001 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf1_), .B(_9269_), .C(_9270_), .Y(_9273_) );
NAND3X1 NAND3X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .B(_9261_), .C(_9266_), .Y(_9274_) );
NAND3X1 NAND3X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_12551_), .B(_9273_), .C(_9274_), .Y(_9275_) );
NAND3X1 NAND3X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_9235_), .B(_9272_), .C(_9275_), .Y(_9276_) );
NAND2X1 NAND2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_12558_), .B(_12560_), .Y(_9277_) );
NAND3X1 NAND3X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_12551_), .B(_9267_), .C(_9271_), .Y(_9278_) );
NAND3X1 NAND3X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_12545_), .B(_9273_), .C(_9274_), .Y(_9279_) );
NAND3X1 NAND3X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_9278_), .B(_9279_), .C(_9277_), .Y(_9280_) );
XNOR2X1 XNOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_11509_), .B(_9102_), .Y(_9281_) );
INVX1 INVX1_1308 ( .gnd(gnd), .vdd(vdd), .A(_9281_), .Y(_9282_) );
NAND3X1 NAND3X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_9276_), .B(_9282_), .C(_9280_), .Y(_9283_) );
AOI21X1 AOI21X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_9278_), .B(_9279_), .C(_9277_), .Y(_9284_) );
AOI21X1 AOI21X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_9272_), .B(_9275_), .C(_9235_), .Y(_9285_) );
OAI21X1 OAI21X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_9285_), .C(_9281_), .Y(_9286_) );
NAND3X1 NAND3X1_2009 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf3_), .B(_9283_), .C(_9286_), .Y(_9287_) );
INVX1 INVX1_1309 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf2_), .Y(_9288_) );
NAND3X1 NAND3X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_9276_), .B(_9281_), .C(_9280_), .Y(_9289_) );
OAI21X1 OAI21X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_9285_), .C(_9282_), .Y(_9290_) );
NAND3X1 NAND3X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_9288_), .B(_9289_), .C(_9290_), .Y(_9291_) );
NAND3X1 NAND3X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_12571_), .B(_9287_), .C(_9291_), .Y(_9292_) );
NAND3X1 NAND3X1_2013 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf1_), .B(_9289_), .C(_9290_), .Y(_9293_) );
NAND3X1 NAND3X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_9288_), .B(_9283_), .C(_9286_), .Y(_9294_) );
NAND3X1 NAND3X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_12577_), .B(_9293_), .C(_9294_), .Y(_9295_) );
NAND3X1 NAND3X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .B(_9295_), .C(_9233_), .Y(_9296_) );
INVX1 INVX1_1310 ( .gnd(gnd), .vdd(vdd), .A(_12583_), .Y(_9297_) );
OAI21X1 OAI21X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_9297_), .B(_12512_), .C(_12582_), .Y(_9298_) );
NAND3X1 NAND3X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_12577_), .B(_9287_), .C(_9291_), .Y(_9299_) );
NAND3X1 NAND3X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_12571_), .B(_9293_), .C(_9294_), .Y(_9300_) );
NAND3X1 NAND3X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_9299_), .B(_9298_), .C(_9300_), .Y(_9301_) );
NAND2X1 NAND2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_9107_), .B(_9109_), .Y(_9302_) );
XNOR2X1 XNOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_11564_), .B(_9302_), .Y(_9303_) );
INVX1 INVX1_1311 ( .gnd(gnd), .vdd(vdd), .A(_9303_), .Y(_9304_) );
NAND3X1 NAND3X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .B(_9301_), .C(_9296_), .Y(_9305_) );
AOI21X1 AOI21X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_9299_), .B(_9300_), .C(_9298_), .Y(_9306_) );
AOI21X1 AOI21X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .B(_9295_), .C(_9233_), .Y(_9307_) );
OAI21X1 OAI21X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_9306_), .B(_9307_), .C(_9303_), .Y(_9308_) );
NAND3X1 NAND3X1_2021 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf1_), .B(_9305_), .C(_9308_), .Y(_9309_) );
INVX1 INVX1_1312 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf0_), .Y(_9310_) );
NAND3X1 NAND3X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_9303_), .B(_9301_), .C(_9296_), .Y(_9311_) );
OAI21X1 OAI21X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_9306_), .B(_9307_), .C(_9304_), .Y(_9312_) );
NAND3X1 NAND3X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_9310_), .B(_9311_), .C(_9312_), .Y(_9313_) );
NAND3X1 NAND3X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_8786_), .B(_9309_), .C(_9313_), .Y(_9314_) );
NAND3X1 NAND3X1_2025 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf3_), .B(_9311_), .C(_9312_), .Y(_9315_) );
NAND3X1 NAND3X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_9310_), .B(_9305_), .C(_9308_), .Y(_9316_) );
NAND3X1 NAND3X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_8792_), .B(_9315_), .C(_9316_), .Y(_9317_) );
NAND3X1 NAND3X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_9231_), .B(_9314_), .C(_9317_), .Y(_9318_) );
NOR3X1 NOR3X1_270 ( .gnd(gnd), .vdd(vdd), .A(_8786_), .B(_12329_), .C(_8790_), .Y(_9319_) );
OAI21X1 OAI21X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_12510_), .C(_8797_), .Y(_9320_) );
NAND3X1 NAND3X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_8792_), .B(_9309_), .C(_9313_), .Y(_9321_) );
NAND3X1 NAND3X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_8786_), .B(_9315_), .C(_9316_), .Y(_9322_) );
NAND3X1 NAND3X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(_9321_), .C(_9322_), .Y(_9323_) );
XNOR2X1 XNOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_11641_), .B(_9116_), .Y(_9324_) );
NAND3X1 NAND3X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_9324_), .B(_9318_), .C(_9323_), .Y(_9325_) );
AOI21X1 AOI21X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .B(_9322_), .C(_9320_), .Y(_9326_) );
AOI21X1 AOI21X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_9314_), .B(_9317_), .C(_9231_), .Y(_9327_) );
INVX1 INVX1_1313 ( .gnd(gnd), .vdd(vdd), .A(_9324_), .Y(_9328_) );
OAI21X1 OAI21X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_9326_), .B(_9327_), .C(_9328_), .Y(_9329_) );
NAND3X1 NAND3X1_2033 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf1_), .B(_9325_), .C(_9329_), .Y(_9330_) );
INVX1 INVX1_1314 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf0_), .Y(_9331_) );
NAND3X1 NAND3X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_9328_), .B(_9318_), .C(_9323_), .Y(_9332_) );
OAI21X1 OAI21X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_9326_), .B(_9327_), .C(_9324_), .Y(_9333_) );
NAND3X1 NAND3X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_9331_), .B(_9332_), .C(_9333_), .Y(_9334_) );
NAND3X1 NAND3X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_8810_), .B(_9330_), .C(_9334_), .Y(_9335_) );
NAND3X1 NAND3X1_2037 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf3_), .B(_9332_), .C(_9333_), .Y(_9336_) );
NAND3X1 NAND3X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_9331_), .B(_9325_), .C(_9329_), .Y(_9337_) );
NAND3X1 NAND3X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_8817_), .B(_9336_), .C(_9337_), .Y(_9338_) );
NAND3X1 NAND3X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_9335_), .C(_9338_), .Y(_9339_) );
NOR3X1 NOR3X1_271 ( .gnd(gnd), .vdd(vdd), .A(_8810_), .B(_8816_), .C(_8814_), .Y(_9340_) );
OAI21X1 OAI21X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_9340_), .B(_12505_), .C(_8822_), .Y(_9341_) );
NAND3X1 NAND3X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_8817_), .B(_9330_), .C(_9334_), .Y(_9342_) );
NAND3X1 NAND3X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_8810_), .B(_9336_), .C(_9337_), .Y(_9343_) );
NAND3X1 NAND3X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_9342_), .B(_9343_), .C(_9341_), .Y(_9344_) );
XNOR2X1 XNOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_11707_), .B(_9124_), .Y(_9345_) );
INVX1 INVX1_1315 ( .gnd(gnd), .vdd(vdd), .A(_9345_), .Y(_9346_) );
NAND3X1 NAND3X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_9346_), .B(_9339_), .C(_9344_), .Y(_9347_) );
AOI21X1 AOI21X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_9342_), .B(_9343_), .C(_9341_), .Y(_9348_) );
AOI21X1 AOI21X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_9335_), .B(_9338_), .C(_9229_), .Y(_9349_) );
OAI21X1 OAI21X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_9348_), .B(_9349_), .C(_9345_), .Y(_9350_) );
NAND3X1 NAND3X1_2045 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf1_), .B(_9347_), .C(_9350_), .Y(_9351_) );
INVX1 INVX1_1316 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf0_), .Y(_9352_) );
NAND3X1 NAND3X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_9345_), .B(_9339_), .C(_9344_), .Y(_9353_) );
OAI21X1 OAI21X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_9348_), .B(_9349_), .C(_9346_), .Y(_9354_) );
NAND3X1 NAND3X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_9352_), .B(_9353_), .C(_9354_), .Y(_9355_) );
NAND3X1 NAND3X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_9351_), .C(_9355_), .Y(_9356_) );
NAND3X1 NAND3X1_2049 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf3_), .B(_9353_), .C(_9354_), .Y(_9357_) );
NAND3X1 NAND3X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_9352_), .B(_9347_), .C(_9350_), .Y(_9358_) );
NAND3X1 NAND3X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_8835_), .B(_9357_), .C(_9358_), .Y(_9359_) );
AOI21X1 AOI21X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_9356_), .B(_9359_), .C(_9227_), .Y(_9360_) );
AOI21X1 AOI21X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_8842_), .C(_12504_), .Y(_9361_) );
AOI21X1 AOI21X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .B(_8849_), .C(_9361_), .Y(_9362_) );
NAND3X1 NAND3X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_8835_), .B(_9351_), .C(_9355_), .Y(_9363_) );
NAND3X1 NAND3X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_9357_), .C(_9358_), .Y(_9364_) );
AOI21X1 AOI21X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_9363_), .B(_9364_), .C(_9362_), .Y(_9365_) );
XNOR2X1 XNOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_11751_), .B(_9132_), .Y(_9366_) );
NOR3X1 NOR3X1_272 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_9366_), .C(_9360_), .Y(_9367_) );
NAND3X1 NAND3X1_2054 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_9363_), .C(_9364_), .Y(_9368_) );
NAND3X1 NAND3X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_9356_), .B(_9359_), .C(_9227_), .Y(_9369_) );
INVX1 INVX1_1317 ( .gnd(gnd), .vdd(vdd), .A(_9366_), .Y(_9370_) );
AOI21X1 AOI21X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_9368_), .B(_9369_), .C(_9370_), .Y(_9371_) );
OAI21X1 OAI21X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_9371_), .C(bloque_datos_85_bF_buf0_), .Y(_9372_) );
INVX1 INVX1_1318 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf4_), .Y(_9373_) );
NAND3X1 NAND3X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_9370_), .B(_9368_), .C(_9369_), .Y(_9374_) );
OAI21X1 OAI21X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_9360_), .B(_9365_), .C(_9366_), .Y(_9375_) );
NAND3X1 NAND3X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_9374_), .C(_9375_), .Y(_9376_) );
NAND3X1 NAND3X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .B(_9376_), .C(_9372_), .Y(_9377_) );
NAND3X1 NAND3X1_2059 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf3_), .B(_9374_), .C(_9375_), .Y(_9378_) );
OAI21X1 OAI21X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_9371_), .C(_9373_), .Y(_9379_) );
NAND3X1 NAND3X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_8867_), .B(_9378_), .C(_9379_), .Y(_9380_) );
NAND3X1 NAND3X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_9225_), .B(_9377_), .C(_9380_), .Y(_9381_) );
NOR3X1 NOR3X1_273 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .B(_12365_), .C(_8865_), .Y(_9382_) );
OAI21X1 OAI21X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_9382_), .B(_12500_), .C(_8872_), .Y(_9383_) );
NAND3X1 NAND3X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_8867_), .B(_9376_), .C(_9372_), .Y(_9384_) );
NAND3X1 NAND3X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .B(_9378_), .C(_9379_), .Y(_9385_) );
NAND3X1 NAND3X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_9384_), .B(_9385_), .C(_9383_), .Y(_9386_) );
XNOR2X1 XNOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_11849_), .B(_9138_), .Y(_9387_) );
NAND3X1 NAND3X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_9387_), .B(_9381_), .C(_9386_), .Y(_9388_) );
AOI21X1 AOI21X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_9384_), .B(_9385_), .C(_9383_), .Y(_9389_) );
AOI21X1 AOI21X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_9377_), .B(_9380_), .C(_9225_), .Y(_9390_) );
INVX1 INVX1_1319 ( .gnd(gnd), .vdd(vdd), .A(_9387_), .Y(_9391_) );
OAI21X1 OAI21X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_9389_), .B(_9390_), .C(_9391_), .Y(_9392_) );
NAND3X1 NAND3X1_2066 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_133_), .B(_9388_), .C(_9392_), .Y(_9393_) );
INVX1 INVX1_1320 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_133_), .Y(_9394_) );
NAND3X1 NAND3X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_9391_), .B(_9381_), .C(_9386_), .Y(_9395_) );
OAI21X1 OAI21X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_9389_), .B(_9390_), .C(_9387_), .Y(_9396_) );
NAND3X1 NAND3X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_9394_), .B(_9395_), .C(_9396_), .Y(_9397_) );
AOI21X1 AOI21X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_9393_), .B(_9397_), .C(_8885_), .Y(_9398_) );
NAND3X1 NAND3X1_2069 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_133_), .B(_9395_), .C(_9396_), .Y(_9399_) );
NAND3X1 NAND3X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_9394_), .B(_9388_), .C(_9392_), .Y(_9400_) );
AOI21X1 AOI21X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_9399_), .B(_9400_), .C(_8892_), .Y(_9401_) );
OAI21X1 OAI21X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_9398_), .B(_9401_), .C(_9223_), .Y(_9402_) );
OAI21X1 OAI21X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_8905_), .B(_8896_), .C(_8890_), .Y(_9403_) );
AOI21X1 AOI21X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_9393_), .B(_9397_), .C(_8892_), .Y(_9404_) );
AOI21X1 AOI21X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_9399_), .B(_9400_), .C(_8885_), .Y(_9405_) );
OAI21X1 OAI21X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_9405_), .C(_9403_), .Y(_9406_) );
NAND3X1 NAND3X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_9147_), .B(_9402_), .C(_9406_), .Y(_9407_) );
NAND3X1 NAND3X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_8892_), .B(_9399_), .C(_9400_), .Y(_9408_) );
NAND3X1 NAND3X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_8885_), .B(_9393_), .C(_9397_), .Y(_9409_) );
AOI21X1 AOI21X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_9408_), .B(_9409_), .C(_9403_), .Y(_9410_) );
NAND3X1 NAND3X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_8885_), .B(_9399_), .C(_9400_), .Y(_9411_) );
NAND3X1 NAND3X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_8892_), .B(_9393_), .C(_9397_), .Y(_9412_) );
AOI21X1 AOI21X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_9412_), .C(_9223_), .Y(_9413_) );
OAI21X1 OAI21X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_9410_), .B(_9413_), .C(_9145_), .Y(_9414_) );
NAND2X1 NAND2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_9407_), .B(_9414_), .Y(_9415_) );
NAND3X1 NAND3X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_9222_), .B(_11926_), .C(_9415_), .Y(_9416_) );
OAI21X1 OAI21X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_9410_), .B(_9413_), .C(_9147_), .Y(_9417_) );
NAND3X1 NAND3X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_9145_), .B(_9402_), .C(_9406_), .Y(_9418_) );
NAND3X1 NAND3X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_11926_), .B(_9418_), .C(_9417_), .Y(_9419_) );
NAND2X1 NAND2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_149_), .B(_9419_), .Y(_9420_) );
NAND3X1 NAND3X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_9221_), .B(_9416_), .C(_9420_), .Y(_9421_) );
NOR2X1 NOR2X1_749 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_149_), .B(_9419_), .Y(_9422_) );
AOI21X1 AOI21X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_11926_), .B(_9415_), .C(_9222_), .Y(_9423_) );
OAI21X1 OAI21X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_9422_), .B(_9423_), .C(_8918_), .Y(_9424_) );
NAND3X1 NAND3X1_2080 ( .gnd(gnd), .vdd(vdd), .A(_9421_), .B(_9220_), .C(_9424_), .Y(_9425_) );
OAI21X1 OAI21X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_8920_), .B(_12498_), .C(_8923_), .Y(_9426_) );
OAI21X1 OAI21X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_9422_), .B(_9423_), .C(_9221_), .Y(_9427_) );
NAND3X1 NAND3X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_8918_), .B(_9416_), .C(_9420_), .Y(_9428_) );
NAND3X1 NAND3X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_9428_), .B(_9427_), .C(_9426_), .Y(_9429_) );
NAND3X1 NAND3X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_9219_), .B(_9425_), .C(_9429_), .Y(_9430_) );
AOI21X1 AOI21X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_9428_), .B(_9427_), .C(_9426_), .Y(_9431_) );
AOI21X1 AOI21X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_9421_), .B(_9424_), .C(_9220_), .Y(_9432_) );
OAI21X1 OAI21X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_9431_), .B(_9432_), .C(_9153_), .Y(_9433_) );
NAND2X1 NAND2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_9430_), .B(_9433_), .Y(_9434_) );
NAND3X1 NAND3X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_9218_), .B(_12010_), .C(_9434_), .Y(_9435_) );
OAI21X1 OAI21X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_9431_), .B(_9432_), .C(_9219_), .Y(_9436_) );
NAND3X1 NAND3X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_9153_), .B(_9425_), .C(_9429_), .Y(_9437_) );
NAND3X1 NAND3X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_12010_), .B(_9437_), .C(_9436_), .Y(_9438_) );
NAND2X1 NAND2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_165_), .B(_9438_), .Y(_9439_) );
NAND3X1 NAND3X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_9217_), .B(_9435_), .C(_9439_), .Y(_9440_) );
NOR2X1 NOR2X1_750 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_165_), .B(_9438_), .Y(_9441_) );
AOI21X1 AOI21X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_12010_), .B(_9434_), .C(_9218_), .Y(_9442_) );
OAI21X1 OAI21X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_9441_), .B(_9442_), .C(_8944_), .Y(_9443_) );
NAND3X1 NAND3X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_9216_), .B(_9440_), .C(_9443_), .Y(_9444_) );
OAI21X1 OAI21X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_12497_), .B(_8946_), .C(_8948_), .Y(_9445_) );
OAI21X1 OAI21X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_9441_), .B(_9442_), .C(_9217_), .Y(_9446_) );
NAND3X1 NAND3X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_9435_), .C(_9439_), .Y(_9447_) );
NAND3X1 NAND3X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_9447_), .B(_9445_), .C(_9446_), .Y(_9448_) );
NAND3X1 NAND3X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .B(_9444_), .C(_9448_), .Y(_9449_) );
NAND2X1 NAND2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_9444_), .B(_9448_), .Y(_9450_) );
AOI21X1 AOI21X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_9162_), .B(_9450_), .C(_12019_), .Y(_9451_) );
NAND3X1 NAND3X1_2092 ( .gnd(gnd), .vdd(vdd), .A(_9215_), .B(_9449_), .C(_9451_), .Y(_9452_) );
AOI21X1 AOI21X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_9447_), .B(_9446_), .C(_9445_), .Y(_9453_) );
AOI21X1 AOI21X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_9440_), .B(_9443_), .C(_9216_), .Y(_9454_) );
OAI21X1 OAI21X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_9453_), .B(_9454_), .C(_9162_), .Y(_9455_) );
NAND3X1 NAND3X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_12018_), .B(_9449_), .C(_9455_), .Y(_9456_) );
NAND2X1 NAND2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_181_), .B(_9456_), .Y(_9457_) );
NAND3X1 NAND3X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_9214_), .B(_9452_), .C(_9457_), .Y(_9458_) );
NOR2X1 NOR2X1_751 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_181_), .B(_9456_), .Y(_9459_) );
AOI21X1 AOI21X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_9449_), .B(_9451_), .C(_9215_), .Y(_9460_) );
OAI21X1 OAI21X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_9460_), .C(_8962_), .Y(_9461_) );
NAND3X1 NAND3X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_9213_), .B(_9458_), .C(_9461_), .Y(_9462_) );
OAI21X1 OAI21X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_8964_), .B(_12494_), .C(_8967_), .Y(_9463_) );
OAI21X1 OAI21X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_9460_), .C(_9214_), .Y(_9464_) );
NAND3X1 NAND3X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_8962_), .B(_9452_), .C(_9457_), .Y(_9465_) );
NAND3X1 NAND3X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_9465_), .B(_9463_), .C(_9464_), .Y(_9466_) );
NAND3X1 NAND3X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_9170_), .B(_9462_), .C(_9466_), .Y(_9467_) );
AOI21X1 AOI21X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_9465_), .B(_9464_), .C(_9463_), .Y(_9468_) );
AOI21X1 AOI21X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_9458_), .B(_9461_), .C(_9213_), .Y(_9469_) );
OAI21X1 OAI21X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_9468_), .B(_9469_), .C(_9169_), .Y(_9470_) );
NAND2X1 NAND2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_9467_), .B(_9470_), .Y(_9471_) );
NAND3X1 NAND3X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_9212_), .B(_12027_), .C(_9471_), .Y(_9472_) );
OAI21X1 OAI21X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_9468_), .B(_9469_), .C(_9170_), .Y(_9473_) );
NAND3X1 NAND3X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_9169_), .B(_9462_), .C(_9466_), .Y(_9474_) );
NAND3X1 NAND3X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_12027_), .B(_9474_), .C(_9473_), .Y(_9475_) );
NAND2X1 NAND2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_197_), .B(_9475_), .Y(_9476_) );
NAND3X1 NAND3X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_9211_), .B(_9472_), .C(_9476_), .Y(_9477_) );
NOR2X1 NOR2X1_752 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_197_), .B(_9475_), .Y(_9478_) );
AOI21X1 AOI21X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_12027_), .B(_9471_), .C(_9212_), .Y(_9479_) );
OAI21X1 OAI21X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_9479_), .C(_8988_), .Y(_9480_) );
NAND3X1 NAND3X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_9477_), .B(_9210_), .C(_9480_), .Y(_9481_) );
OAI21X1 OAI21X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_8990_), .B(_12492_), .C(_8993_), .Y(_9482_) );
OAI21X1 OAI21X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_9479_), .C(_9211_), .Y(_9483_) );
NAND3X1 NAND3X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_8988_), .B(_9472_), .C(_9476_), .Y(_9484_) );
NAND3X1 NAND3X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9483_), .C(_9482_), .Y(_9485_) );
NAND3X1 NAND3X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_9178_), .B(_9481_), .C(_9485_), .Y(_9486_) );
AOI21X1 AOI21X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9483_), .C(_9482_), .Y(_9487_) );
AOI21X1 AOI21X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_9477_), .B(_9480_), .C(_9210_), .Y(_9488_) );
OAI21X1 OAI21X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_9487_), .B(_9488_), .C(_9177_), .Y(_9489_) );
NAND2X1 NAND2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_9486_), .B(_9489_), .Y(_9490_) );
NAND3X1 NAND3X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_9209_), .B(_12035_), .C(_9490_), .Y(_9491_) );
OAI21X1 OAI21X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_9487_), .B(_9488_), .C(_9178_), .Y(_9492_) );
NAND3X1 NAND3X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_9177_), .B(_9481_), .C(_9485_), .Y(_9493_) );
NAND3X1 NAND3X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_12035_), .B(_9493_), .C(_9492_), .Y(_9494_) );
NAND2X1 NAND2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_213_), .B(_9494_), .Y(_9495_) );
NAND3X1 NAND3X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_9491_), .C(_9495_), .Y(_9496_) );
NOR2X1 NOR2X1_753 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_213_), .B(_9494_), .Y(_9497_) );
AOI21X1 AOI21X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_12035_), .B(_9490_), .C(_9209_), .Y(_9498_) );
OAI21X1 OAI21X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_9497_), .B(_9498_), .C(_9009_), .Y(_9499_) );
NAND3X1 NAND3X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_9496_), .B(_9207_), .C(_9499_), .Y(_9500_) );
OAI21X1 OAI21X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_9011_), .B(_12490_), .C(_9015_), .Y(_9501_) );
OAI21X1 OAI21X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_9497_), .B(_9498_), .C(_9208_), .Y(_9502_) );
NAND3X1 NAND3X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_9009_), .B(_9491_), .C(_9495_), .Y(_9503_) );
NAND3X1 NAND3X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_9503_), .B(_9501_), .C(_9502_), .Y(_9504_) );
NAND3X1 NAND3X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_9186_), .B(_9500_), .C(_9504_), .Y(_9505_) );
AOI21X1 AOI21X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_9503_), .B(_9502_), .C(_9501_), .Y(_9506_) );
AOI21X1 AOI21X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_9496_), .B(_9499_), .C(_9207_), .Y(_9507_) );
OAI21X1 OAI21X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_9506_), .B(_9507_), .C(_9185_), .Y(_9508_) );
NAND2X1 NAND2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_9505_), .B(_9508_), .Y(_9509_) );
NAND3X1 NAND3X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_9206_), .B(_12044_), .C(_9509_), .Y(_9510_) );
OAI21X1 OAI21X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_9506_), .B(_9507_), .C(_9186_), .Y(_9511_) );
NAND3X1 NAND3X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_9500_), .C(_9504_), .Y(_9512_) );
NAND3X1 NAND3X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_12044_), .B(_9512_), .C(_9511_), .Y(_9513_) );
NAND2X1 NAND2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_229_), .B(_9513_), .Y(_9514_) );
NAND3X1 NAND3X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_9205_), .B(_9510_), .C(_9514_), .Y(_9515_) );
NOR2X1 NOR2X1_754 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_229_), .B(_9513_), .Y(_9516_) );
AOI21X1 AOI21X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_12044_), .B(_9509_), .C(_9206_), .Y(_9517_) );
OAI21X1 OAI21X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_9516_), .B(_9517_), .C(_9036_), .Y(_9518_) );
NAND3X1 NAND3X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_9204_), .B(_9515_), .C(_9518_), .Y(_9519_) );
OAI21X1 OAI21X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_12488_), .B(_9038_), .C(_9041_), .Y(_9520_) );
OAI21X1 OAI21X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_9516_), .B(_9517_), .C(_9205_), .Y(_9521_) );
NAND3X1 NAND3X1_2120 ( .gnd(gnd), .vdd(vdd), .A(_9036_), .B(_9510_), .C(_9514_), .Y(_9522_) );
NAND3X1 NAND3X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_9520_), .B(_9522_), .C(_9521_), .Y(_9523_) );
NAND3X1 NAND3X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_9193_), .B(_9519_), .C(_9523_), .Y(_9524_) );
NAND2X1 NAND2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_9519_), .B(_9523_), .Y(_9525_) );
AOI21X1 AOI21X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(_9525_), .C(_12241_), .Y(_9526_) );
NAND3X1 NAND3X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(_9524_), .C(_9526_), .Y(_9527_) );
AOI21X1 AOI21X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_9522_), .B(_9521_), .C(_9520_), .Y(_9528_) );
AOI21X1 AOI21X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_9515_), .B(_9518_), .C(_9204_), .Y(_9529_) );
OAI21X1 OAI21X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_9528_), .B(_9529_), .C(_9194_), .Y(_9530_) );
NAND3X1 NAND3X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_12052_), .B(_9524_), .C(_9530_), .Y(_9531_) );
NAND2X1 NAND2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_245_), .B(_9531_), .Y(_9532_) );
NAND3X1 NAND3X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_9053_), .B(_9527_), .C(_9532_), .Y(_9533_) );
INVX1 INVX1_1321 ( .gnd(gnd), .vdd(vdd), .A(_9053_), .Y(_9534_) );
NOR2X1 NOR2X1_755 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_245_), .B(_9531_), .Y(_9535_) );
AOI21X1 AOI21X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_9524_), .B(_9526_), .C(_9203_), .Y(_9536_) );
OAI21X1 OAI21X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_9535_), .B(_9536_), .C(_9534_), .Y(_9537_) );
NAND3X1 NAND3X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_9533_), .B(_9202_), .C(_9537_), .Y(_9538_) );
AOI21X1 AOI21X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_12486_), .C(_9065_), .Y(_9539_) );
NOR3X1 NOR3X1_274 ( .gnd(gnd), .vdd(vdd), .A(_9534_), .B(_9536_), .C(_9535_), .Y(_9540_) );
AOI21X1 AOI21X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_9527_), .B(_9532_), .C(_9053_), .Y(_9541_) );
OAI21X1 OAI21X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_9540_), .B(_9541_), .C(_9539_), .Y(_9542_) );
NAND3X1 NAND3X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_9201_), .B(_9538_), .C(_9542_), .Y(_9543_) );
INVX1 INVX1_1322 ( .gnd(gnd), .vdd(vdd), .A(_9201_), .Y(_9544_) );
NAND3X1 NAND3X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_9533_), .B(_9539_), .C(_9537_), .Y(_9545_) );
OAI21X1 OAI21X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_9540_), .B(_9541_), .C(_9202_), .Y(_9546_) );
NAND3X1 NAND3X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_9544_), .B(_9545_), .C(_9546_), .Y(_9547_) );
NAND2X1 NAND2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_9543_), .B(_9547_), .Y(_9548_) );
XNOR2X1 XNOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_9548_), .B(_9077_), .Y(module_2_H_5_) );
AOI21X1 AOI21X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_9543_), .B(_9547_), .C(_9077_), .Y(_9549_) );
AOI21X1 AOI21X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_9533_), .B(_9202_), .C(_9541_), .Y(_9550_) );
AOI21X1 AOI21X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_9510_), .B(_9514_), .C(_9036_), .Y(_9551_) );
AOI21X1 AOI21X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_9522_), .B(_9520_), .C(_9551_), .Y(_9552_) );
INVX1 INVX1_1323 ( .gnd(gnd), .vdd(vdd), .A(_12222_), .Y(_9553_) );
INVX1 INVX1_1324 ( .gnd(gnd), .vdd(vdd), .A(_12223_), .Y(_9554_) );
NOR2X1 NOR2X1_756 ( .gnd(gnd), .vdd(vdd), .A(_9554_), .B(_9553_), .Y(_9555_) );
INVX1 INVX1_1325 ( .gnd(gnd), .vdd(vdd), .A(_9555_), .Y(_9556_) );
AOI21X1 AOI21X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_9491_), .B(_9495_), .C(_9009_), .Y(_9557_) );
AOI21X1 AOI21X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_9503_), .B(_9501_), .C(_9557_), .Y(_9558_) );
INVX1 INVX1_1326 ( .gnd(gnd), .vdd(vdd), .A(_12212_), .Y(_9559_) );
AOI21X1 AOI21X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_9472_), .B(_9476_), .C(_8988_), .Y(_9560_) );
AOI21X1 AOI21X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(_9560_), .Y(_9561_) );
NOR2X1 NOR2X1_757 ( .gnd(gnd), .vdd(vdd), .A(_12202_), .B(_12201_), .Y(_9562_) );
INVX2 INVX2_332 ( .gnd(gnd), .vdd(vdd), .A(_9562_), .Y(_9563_) );
NOR3X1 NOR3X1_275 ( .gnd(gnd), .vdd(vdd), .A(_9214_), .B(_9460_), .C(_9459_), .Y(_9564_) );
OAI21X1 OAI21X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_9564_), .B(_9213_), .C(_9464_), .Y(_9565_) );
INVX2 INVX2_333 ( .gnd(gnd), .vdd(vdd), .A(_12194_), .Y(_9566_) );
AOI21X1 AOI21X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_9435_), .B(_9439_), .C(_8944_), .Y(_9567_) );
AOI21X1 AOI21X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_9447_), .B(_9445_), .C(_9567_), .Y(_9568_) );
INVX1 INVX1_1327 ( .gnd(gnd), .vdd(vdd), .A(_9427_), .Y(_9569_) );
AOI21X1 AOI21X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_9428_), .B(_9426_), .C(_9569_), .Y(_9570_) );
NOR2X1 NOR2X1_758 ( .gnd(gnd), .vdd(vdd), .A(_12173_), .B(_12174_), .Y(_9571_) );
INVX1 INVX1_1328 ( .gnd(gnd), .vdd(vdd), .A(_9571_), .Y(_9572_) );
OAI21X1 OAI21X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_9223_), .C(_9408_), .Y(_9573_) );
INVX2 INVX2_334 ( .gnd(gnd), .vdd(vdd), .A(_9399_), .Y(_9574_) );
AOI21X1 AOI21X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_9372_), .C(_8867_), .Y(_9575_) );
OAI21X1 OAI21X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_9575_), .B(_9225_), .C(_9384_), .Y(_9576_) );
INVX2 INVX2_335 ( .gnd(gnd), .vdd(vdd), .A(_9372_), .Y(_9577_) );
NAND2X1 NAND2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_9356_), .B(_9369_), .Y(_9578_) );
INVX2 INVX2_336 ( .gnd(gnd), .vdd(vdd), .A(_9351_), .Y(_9579_) );
NAND2X1 NAND2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_9342_), .B(_9344_), .Y(_9580_) );
INVX2 INVX2_337 ( .gnd(gnd), .vdd(vdd), .A(_9330_), .Y(_9581_) );
NAND2X1 NAND2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .B(_9323_), .Y(_9582_) );
INVX2 INVX2_338 ( .gnd(gnd), .vdd(vdd), .A(_9309_), .Y(_9583_) );
NAND2X1 NAND2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_9299_), .B(_9301_), .Y(_9584_) );
INVX2 INVX2_339 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .Y(_9585_) );
INVX1 INVX1_1329 ( .gnd(gnd), .vdd(vdd), .A(_9279_), .Y(_9586_) );
OAI21X1 OAI21X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_9586_), .B(_9235_), .C(_9278_), .Y(_9587_) );
INVX2 INVX2_340 ( .gnd(gnd), .vdd(vdd), .A(_9267_), .Y(_9588_) );
NAND3X1 NAND3X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_12530_), .B(_9247_), .C(_9251_), .Y(_9589_) );
INVX1 INVX1_1330 ( .gnd(gnd), .vdd(vdd), .A(_9247_), .Y(_9590_) );
NAND2X1 NAND2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_12069_), .B(_12073_), .Y(_9591_) );
INVX1 INVX1_1331 ( .gnd(gnd), .vdd(vdd), .A(_9591_), .Y(_9592_) );
INVX1 INVX1_1332 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_6_), .Y(_9593_) );
AND2X2 AND2X2_210 ( .gnd(gnd), .vdd(vdd), .A(_9244_), .B(_9593_), .Y(_9594_) );
NOR2X1 NOR2X1_759 ( .gnd(gnd), .vdd(vdd), .A(_9593_), .B(_9244_), .Y(_9595_) );
OAI21X1 OAI21X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_9594_), .B(_9595_), .C(_9592_), .Y(_9596_) );
NOR2X1 NOR2X1_760 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .B(_9594_), .Y(_9597_) );
OAI21X1 OAI21X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_12070_), .B(_12071_), .C(_9597_), .Y(_9598_) );
NAND3X1 NAND3X1_2131 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_22_), .B(_9596_), .C(_9598_), .Y(_9599_) );
INVX1 INVX1_1333 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_22_), .Y(_9600_) );
OAI21X1 OAI21X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_9594_), .B(_9595_), .C(_9591_), .Y(_9601_) );
NAND2X1 NAND2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_9592_), .B(_9597_), .Y(_9602_) );
NAND3X1 NAND3X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_9600_), .B(_9601_), .C(_9602_), .Y(_9603_) );
NAND3X1 NAND3X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_9590_), .B(_9603_), .C(_9599_), .Y(_9604_) );
AOI21X1 AOI21X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_9601_), .B(_9602_), .C(_9600_), .Y(_9605_) );
AOI21X1 AOI21X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_9596_), .B(_9598_), .C(module_2_W_22_), .Y(_9606_) );
OAI21X1 OAI21X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_9606_), .B(_9605_), .C(_9247_), .Y(_9607_) );
NAND2X1 NAND2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_9604_), .B(_9607_), .Y(_9608_) );
AOI21X1 AOI21X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_9589_), .B(_9259_), .C(_9608_), .Y(_9609_) );
INVX1 INVX1_1334 ( .gnd(gnd), .vdd(vdd), .A(_9609_), .Y(_9610_) );
OAI21X1 OAI21X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_9237_), .B(_9256_), .C(_9589_), .Y(_9611_) );
INVX1 INVX1_1335 ( .gnd(gnd), .vdd(vdd), .A(_9608_), .Y(_9612_) );
OR2X2 OR2X2_233 ( .gnd(gnd), .vdd(vdd), .A(_9612_), .B(_9611_), .Y(_9613_) );
INVX2 INVX2_341 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_10_), .Y(_9614_) );
NOR2X1 NOR2X1_761 ( .gnd(gnd), .vdd(vdd), .A(_12082_), .B(_12080_), .Y(_9615_) );
XNOR2X1 XNOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_9615_), .B(_9614_), .Y(_9616_) );
NAND3X1 NAND3X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_9610_), .B(_9616_), .C(_9613_), .Y(_9617_) );
NOR2X1 NOR2X1_762 ( .gnd(gnd), .vdd(vdd), .A(_9611_), .B(_9612_), .Y(_9618_) );
INVX1 INVX1_1336 ( .gnd(gnd), .vdd(vdd), .A(_9616_), .Y(_9619_) );
OAI21X1 OAI21X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_9618_), .B(_9609_), .C(_9619_), .Y(_9620_) );
NAND3X1 NAND3X1_2135 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf3_), .B(_9620_), .C(_9617_), .Y(_9621_) );
INVX2 INVX2_342 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf2_), .Y(_9622_) );
NAND3X1 NAND3X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_9610_), .B(_9619_), .C(_9613_), .Y(_9623_) );
OAI21X1 OAI21X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_9618_), .B(_9609_), .C(_9616_), .Y(_9624_) );
NAND3X1 NAND3X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_9622_), .B(_9624_), .C(_9623_), .Y(_9625_) );
NAND3X1 NAND3X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_9588_), .B(_9621_), .C(_9625_), .Y(_9626_) );
NAND3X1 NAND3X1_2139 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf1_), .B(_9624_), .C(_9623_), .Y(_9627_) );
NAND3X1 NAND3X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_9622_), .B(_9620_), .C(_9617_), .Y(_9628_) );
NAND3X1 NAND3X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_9267_), .B(_9627_), .C(_9628_), .Y(_9629_) );
NAND3X1 NAND3X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_9587_), .B(_9626_), .C(_9629_), .Y(_9630_) );
INVX1 INVX1_1337 ( .gnd(gnd), .vdd(vdd), .A(_9278_), .Y(_9631_) );
NOR2X1 NOR2X1_763 ( .gnd(gnd), .vdd(vdd), .A(_9631_), .B(_9285_), .Y(_9632_) );
AOI21X1 AOI21X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_9627_), .B(_9628_), .C(_9267_), .Y(_9633_) );
AOI21X1 AOI21X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_9621_), .B(_9625_), .C(_9588_), .Y(_9634_) );
OAI21X1 OAI21X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_9633_), .B(_9634_), .C(_9632_), .Y(_9635_) );
NOR2X1 NOR2X1_764 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_12099_), .Y(_9636_) );
NAND2X1 NAND2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_26_), .B(module_2_W_10_), .Y(_9637_) );
INVX1 INVX1_1338 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_26_), .Y(_9638_) );
NAND2X1 NAND2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_9638_), .B(_9614_), .Y(_9639_) );
AND2X2 AND2X2_211 ( .gnd(gnd), .vdd(vdd), .A(_9639_), .B(_9637_), .Y(_9640_) );
NAND2X1 NAND2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_9640_), .Y(_9641_) );
NAND2X1 NAND2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_9637_), .B(_9639_), .Y(_9642_) );
OAI21X1 OAI21X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_9095_), .B(_9096_), .C(_9642_), .Y(_9643_) );
NAND3X1 NAND3X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_9641_), .B(_9643_), .C(_9101_), .Y(_9644_) );
OAI21X1 OAI21X1_1501 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_24_), .B(module_2_W_8_), .C(_9099_), .Y(_9645_) );
INVX1 INVX1_1339 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .Y(_9646_) );
NOR2X1 NOR2X1_765 ( .gnd(gnd), .vdd(vdd), .A(_9646_), .B(_9642_), .Y(_9647_) );
NOR2X1 NOR2X1_766 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_9640_), .Y(_9648_) );
OAI21X1 OAI21X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_9648_), .B(_9647_), .C(_9645_), .Y(_9649_) );
NAND2X1 NAND2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_9649_), .B(_9644_), .Y(_9650_) );
XNOR2X1 XNOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_9636_), .B(_9650_), .Y(_9651_) );
NAND3X1 NAND3X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_9630_), .B(_9651_), .C(_9635_), .Y(_9652_) );
NAND3X1 NAND3X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_9267_), .B(_9621_), .C(_9625_), .Y(_9653_) );
NAND3X1 NAND3X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_9588_), .B(_9627_), .C(_9628_), .Y(_9654_) );
AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_9278_), .B(_9280_), .C(_9653_), .D(_9654_), .Y(_9655_) );
AOI21X1 AOI21X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_9626_), .B(_9629_), .C(_9587_), .Y(_9656_) );
INVX1 INVX1_1340 ( .gnd(gnd), .vdd(vdd), .A(_9651_), .Y(_9657_) );
OAI21X1 OAI21X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_9655_), .B(_9656_), .C(_9657_), .Y(_9658_) );
NAND3X1 NAND3X1_2147 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf3_), .B(_9652_), .C(_9658_), .Y(_9659_) );
INVX1 INVX1_1341 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf2_), .Y(_9660_) );
NAND3X1 NAND3X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_9630_), .B(_9657_), .C(_9635_), .Y(_9661_) );
OAI21X1 OAI21X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_9655_), .B(_9656_), .C(_9651_), .Y(_9662_) );
NAND3X1 NAND3X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_9660_), .B(_9661_), .C(_9662_), .Y(_9663_) );
NAND3X1 NAND3X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_9585_), .B(_9659_), .C(_9663_), .Y(_9664_) );
NAND3X1 NAND3X1_2151 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf1_), .B(_9661_), .C(_9662_), .Y(_9665_) );
NAND3X1 NAND3X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_9660_), .B(_9652_), .C(_9658_), .Y(_9666_) );
NAND3X1 NAND3X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .B(_9665_), .C(_9666_), .Y(_9667_) );
NAND3X1 NAND3X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_9664_), .B(_9667_), .C(_9584_), .Y(_9668_) );
AND2X2 AND2X2_212 ( .gnd(gnd), .vdd(vdd), .A(_9301_), .B(_9299_), .Y(_9669_) );
AOI21X1 AOI21X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_9665_), .B(_9666_), .C(_9287_), .Y(_9670_) );
AOI21X1 AOI21X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_9659_), .B(_9663_), .C(_9585_), .Y(_9671_) );
OAI21X1 OAI21X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_9670_), .B(_9671_), .C(_9669_), .Y(_9672_) );
NOR2X1 NOR2X1_767 ( .gnd(gnd), .vdd(vdd), .A(_12109_), .B(_12106_), .Y(_9673_) );
NOR2X1 NOR2X1_768 ( .gnd(gnd), .vdd(vdd), .A(_9094_), .B(_9108_), .Y(_9674_) );
INVX1 INVX1_1342 ( .gnd(gnd), .vdd(vdd), .A(_9106_), .Y(_9675_) );
INVX1 INVX1_1343 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .Y(_9676_) );
NAND2X1 NAND2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_9676_), .B(_9650_), .Y(_9677_) );
NAND3X1 NAND3X1_2155 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .B(_9649_), .C(_9644_), .Y(_9678_) );
NAND2X1 NAND2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_9678_), .B(_9677_), .Y(_9679_) );
NOR2X1 NOR2X1_769 ( .gnd(gnd), .vdd(vdd), .A(_9675_), .B(_9679_), .Y(_9680_) );
AOI21X1 AOI21X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_9678_), .B(_9677_), .C(_9106_), .Y(_9681_) );
NOR2X1 NOR2X1_770 ( .gnd(gnd), .vdd(vdd), .A(_9681_), .B(_9680_), .Y(_9682_) );
NAND2X1 NAND2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_9674_), .B(_9682_), .Y(_9683_) );
OAI21X1 OAI21X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_9680_), .B(_9681_), .C(_9109_), .Y(_9684_) );
NAND2X1 NAND2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_9684_), .B(_9683_), .Y(_9685_) );
XNOR2X1 XNOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_9673_), .B(_9685_), .Y(_9686_) );
NAND3X1 NAND3X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_9668_), .B(_9686_), .C(_9672_), .Y(_9687_) );
NAND3X1 NAND3X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .B(_9659_), .C(_9663_), .Y(_9688_) );
NAND3X1 NAND3X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_9585_), .B(_9665_), .C(_9666_), .Y(_9689_) );
AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_9299_), .B(_9301_), .C(_9688_), .D(_9689_), .Y(_9690_) );
AOI21X1 AOI21X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_9664_), .B(_9667_), .C(_9584_), .Y(_9691_) );
INVX1 INVX1_1344 ( .gnd(gnd), .vdd(vdd), .A(_9686_), .Y(_9692_) );
OAI21X1 OAI21X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_9690_), .B(_9691_), .C(_9692_), .Y(_9693_) );
NAND3X1 NAND3X1_2159 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf1_), .B(_9693_), .C(_9687_), .Y(_9694_) );
INVX1 INVX1_1345 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf0_), .Y(_9695_) );
NAND3X1 NAND3X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_9668_), .B(_9692_), .C(_9672_), .Y(_9696_) );
OAI21X1 OAI21X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_9690_), .B(_9691_), .C(_9686_), .Y(_9697_) );
NAND3X1 NAND3X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_9695_), .B(_9697_), .C(_9696_), .Y(_9698_) );
NAND3X1 NAND3X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_9583_), .B(_9694_), .C(_9698_), .Y(_9699_) );
NAND3X1 NAND3X1_2163 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf3_), .B(_9697_), .C(_9696_), .Y(_9700_) );
NAND3X1 NAND3X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_9695_), .B(_9693_), .C(_9687_), .Y(_9701_) );
NAND3X1 NAND3X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_9309_), .B(_9700_), .C(_9701_), .Y(_9702_) );
NAND3X1 NAND3X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_9699_), .B(_9702_), .C(_9582_), .Y(_9703_) );
AND2X2 AND2X2_213 ( .gnd(gnd), .vdd(vdd), .A(_9323_), .B(_9321_), .Y(_9704_) );
AOI21X1 AOI21X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_9700_), .B(_9701_), .C(_9309_), .Y(_9705_) );
AOI21X1 AOI21X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_9694_), .B(_9698_), .C(_9583_), .Y(_9706_) );
OAI21X1 OAI21X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_9705_), .B(_9706_), .C(_9704_), .Y(_9707_) );
INVX2 INVX2_343 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf3_), .Y(_9708_) );
AND2X2 AND2X2_214 ( .gnd(gnd), .vdd(vdd), .A(_9682_), .B(_9674_), .Y(_9709_) );
INVX1 INVX1_1346 ( .gnd(gnd), .vdd(vdd), .A(_9684_), .Y(_9710_) );
OAI21X1 OAI21X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_9709_), .B(_9710_), .C(_9708_), .Y(_9711_) );
OR2X2 OR2X2_234 ( .gnd(gnd), .vdd(vdd), .A(_9685_), .B(_9708_), .Y(_9712_) );
NAND3X1 NAND3X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_9711_), .C(_9712_), .Y(_9713_) );
INVX1 INVX1_1347 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .Y(_9714_) );
INVX1 INVX1_1348 ( .gnd(gnd), .vdd(vdd), .A(_9711_), .Y(_9715_) );
NOR2X1 NOR2X1_771 ( .gnd(gnd), .vdd(vdd), .A(_9708_), .B(_9685_), .Y(_9716_) );
OAI21X1 OAI21X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_9715_), .B(_9716_), .C(_9714_), .Y(_9717_) );
NAND2X1 NAND2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_9713_), .B(_9717_), .Y(_9718_) );
OR2X2 OR2X2_235 ( .gnd(gnd), .vdd(vdd), .A(_9718_), .B(_9115_), .Y(_9719_) );
NOR3X1 NOR3X1_276 ( .gnd(gnd), .vdd(vdd), .A(_9714_), .B(_9716_), .C(_9715_), .Y(_9720_) );
AOI21X1 AOI21X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_9711_), .B(_9712_), .C(_9112_), .Y(_9721_) );
OAI21X1 OAI21X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_9720_), .B(_9721_), .C(_9115_), .Y(_9722_) );
NAND2X1 NAND2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_9722_), .B(_9719_), .Y(_9723_) );
XNOR2X1 XNOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_12338_), .B(_9723_), .Y(_9724_) );
NAND3X1 NAND3X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_9703_), .B(_9724_), .C(_9707_), .Y(_9725_) );
NAND3X1 NAND3X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_9309_), .B(_9694_), .C(_9698_), .Y(_9726_) );
NAND3X1 NAND3X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_9583_), .B(_9700_), .C(_9701_), .Y(_9727_) );
AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .B(_9323_), .C(_9726_), .D(_9727_), .Y(_9728_) );
AOI21X1 AOI21X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_9699_), .B(_9702_), .C(_9582_), .Y(_9729_) );
INVX1 INVX1_1349 ( .gnd(gnd), .vdd(vdd), .A(_9724_), .Y(_9730_) );
OAI21X1 OAI21X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_9728_), .B(_9729_), .C(_9730_), .Y(_9731_) );
NAND3X1 NAND3X1_2171 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf1_), .B(_9725_), .C(_9731_), .Y(_9732_) );
INVX1 INVX1_1350 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf0_), .Y(_9733_) );
OAI21X1 OAI21X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_9728_), .B(_9729_), .C(_9724_), .Y(_9734_) );
NAND3X1 NAND3X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_9703_), .B(_9730_), .C(_9707_), .Y(_9735_) );
NAND3X1 NAND3X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_9733_), .B(_9735_), .C(_9734_), .Y(_9736_) );
NAND3X1 NAND3X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_9581_), .B(_9732_), .C(_9736_), .Y(_9737_) );
NAND3X1 NAND3X1_2175 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf3_), .B(_9735_), .C(_9734_), .Y(_9738_) );
NAND3X1 NAND3X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_9733_), .B(_9725_), .C(_9731_), .Y(_9739_) );
NAND3X1 NAND3X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_9330_), .B(_9738_), .C(_9739_), .Y(_9740_) );
NAND3X1 NAND3X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_9737_), .B(_9740_), .C(_9580_), .Y(_9741_) );
AND2X2 AND2X2_215 ( .gnd(gnd), .vdd(vdd), .A(_9344_), .B(_9342_), .Y(_9742_) );
AOI21X1 AOI21X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_9738_), .B(_9739_), .C(_9330_), .Y(_9743_) );
AOI21X1 AOI21X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_9732_), .B(_9736_), .C(_9581_), .Y(_9744_) );
OAI21X1 OAI21X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_9743_), .B(_9744_), .C(_9742_), .Y(_9745_) );
INVX1 INVX1_1351 ( .gnd(gnd), .vdd(vdd), .A(_9120_), .Y(_9746_) );
INVX1 INVX1_1352 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf1_), .Y(_9747_) );
NOR2X1 NOR2X1_772 ( .gnd(gnd), .vdd(vdd), .A(_9115_), .B(_9718_), .Y(_9748_) );
INVX1 INVX1_1353 ( .gnd(gnd), .vdd(vdd), .A(_9722_), .Y(_9749_) );
OAI21X1 OAI21X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_9749_), .B(_9748_), .C(_9747_), .Y(_9750_) );
INVX1 INVX1_1354 ( .gnd(gnd), .vdd(vdd), .A(_9750_), .Y(_9751_) );
NOR2X1 NOR2X1_773 ( .gnd(gnd), .vdd(vdd), .A(_9747_), .B(_9723_), .Y(_9752_) );
NOR3X1 NOR3X1_277 ( .gnd(gnd), .vdd(vdd), .A(_9751_), .B(_9746_), .C(_9752_), .Y(_9753_) );
NOR2X1 NOR2X1_774 ( .gnd(gnd), .vdd(vdd), .A(_9748_), .B(_9749_), .Y(_9754_) );
NAND2X1 NAND2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf0_), .B(_9754_), .Y(_9755_) );
AOI21X1 AOI21X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_9750_), .B(_9755_), .C(_9120_), .Y(_9756_) );
NOR3X1 NOR3X1_278 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_9756_), .C(_9753_), .Y(_9757_) );
INVX2 INVX2_344 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .Y(_9758_) );
NAND3X1 NAND3X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_9120_), .B(_9750_), .C(_9755_), .Y(_9759_) );
OAI21X1 OAI21X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_9752_), .B(_9751_), .C(_9746_), .Y(_9760_) );
AOI21X1 AOI21X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_9759_), .B(_9760_), .C(_9758_), .Y(_9761_) );
NOR2X1 NOR2X1_775 ( .gnd(gnd), .vdd(vdd), .A(_9761_), .B(_9757_), .Y(_9762_) );
OAI21X1 OAI21X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_12129_), .B(_12130_), .C(_9762_), .Y(_9763_) );
NOR2X1 NOR2X1_776 ( .gnd(gnd), .vdd(vdd), .A(_12130_), .B(_12129_), .Y(_9764_) );
OAI21X1 OAI21X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_9757_), .B(_9761_), .C(_9764_), .Y(_9765_) );
NAND2X1 NAND2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_9763_), .B(_9765_), .Y(_9766_) );
NAND3X1 NAND3X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_9741_), .B(_9766_), .C(_9745_), .Y(_9767_) );
NAND3X1 NAND3X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_9330_), .B(_9732_), .C(_9736_), .Y(_9768_) );
NAND3X1 NAND3X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_9581_), .B(_9738_), .C(_9739_), .Y(_9769_) );
AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_9342_), .B(_9344_), .C(_9768_), .D(_9769_), .Y(_9770_) );
AOI21X1 AOI21X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_9737_), .B(_9740_), .C(_9580_), .Y(_9771_) );
INVX1 INVX1_1355 ( .gnd(gnd), .vdd(vdd), .A(_9766_), .Y(_9772_) );
OAI21X1 OAI21X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_9770_), .B(_9771_), .C(_9772_), .Y(_9773_) );
NAND3X1 NAND3X1_2183 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf1_), .B(_9767_), .C(_9773_), .Y(_9774_) );
INVX1 INVX1_1356 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf0_), .Y(_9775_) );
OAI21X1 OAI21X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_9770_), .B(_9771_), .C(_9766_), .Y(_9776_) );
NAND3X1 NAND3X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_9741_), .B(_9772_), .C(_9745_), .Y(_9777_) );
NAND3X1 NAND3X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_9775_), .B(_9777_), .C(_9776_), .Y(_9778_) );
NAND3X1 NAND3X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_9579_), .B(_9774_), .C(_9778_), .Y(_9779_) );
NAND3X1 NAND3X1_2187 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf3_), .B(_9777_), .C(_9776_), .Y(_9780_) );
NAND3X1 NAND3X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_9775_), .B(_9767_), .C(_9773_), .Y(_9781_) );
NAND3X1 NAND3X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_9351_), .B(_9780_), .C(_9781_), .Y(_9782_) );
NAND3X1 NAND3X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_9779_), .B(_9782_), .C(_9578_), .Y(_9783_) );
AND2X2 AND2X2_216 ( .gnd(gnd), .vdd(vdd), .A(_9369_), .B(_9356_), .Y(_9784_) );
AOI21X1 AOI21X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_9780_), .B(_9781_), .C(_9351_), .Y(_9785_) );
AOI21X1 AOI21X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_9774_), .B(_9778_), .C(_9579_), .Y(_9786_) );
OAI21X1 OAI21X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_9785_), .B(_9786_), .C(_9784_), .Y(_9787_) );
INVX1 INVX1_1357 ( .gnd(gnd), .vdd(vdd), .A(_9128_), .Y(_9788_) );
NAND3X1 NAND3X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_9759_), .B(_9760_), .C(_9758_), .Y(_9789_) );
OAI21X1 OAI21X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_9753_), .B(_9756_), .C(_9123_), .Y(_9790_) );
AOI21X1 AOI21X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_9789_), .B(_9790_), .C(bloque_datos_58_bF_buf2_), .Y(_9791_) );
INVX1 INVX1_1358 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf1_), .Y(_9792_) );
NOR3X1 NOR3X1_279 ( .gnd(gnd), .vdd(vdd), .A(_9792_), .B(_9761_), .C(_9757_), .Y(_9793_) );
NOR3X1 NOR3X1_280 ( .gnd(gnd), .vdd(vdd), .A(_9788_), .B(_9791_), .C(_9793_), .Y(_9794_) );
OAI21X1 OAI21X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_9757_), .B(_9761_), .C(_9792_), .Y(_9795_) );
NAND3X1 NAND3X1_2192 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf0_), .B(_9789_), .C(_9790_), .Y(_9796_) );
AOI21X1 AOI21X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_9796_), .B(_9795_), .C(_9128_), .Y(_9797_) );
NOR3X1 NOR3X1_281 ( .gnd(gnd), .vdd(vdd), .A(_9131_), .B(_9797_), .C(_9794_), .Y(_9798_) );
NOR2X1 NOR2X1_777 ( .gnd(gnd), .vdd(vdd), .A(_9091_), .B(_9130_), .Y(_9799_) );
NAND3X1 NAND3X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_9128_), .B(_9796_), .C(_9795_), .Y(_9800_) );
OAI21X1 OAI21X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_9793_), .B(_9791_), .C(_9788_), .Y(_9801_) );
AOI21X1 AOI21X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_9800_), .B(_9801_), .C(_9799_), .Y(_9802_) );
NOR2X1 NOR2X1_778 ( .gnd(gnd), .vdd(vdd), .A(_9802_), .B(_9798_), .Y(_9803_) );
OAI21X1 OAI21X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_12149_), .B(_12150_), .C(_9803_), .Y(_9804_) );
NOR2X1 NOR2X1_779 ( .gnd(gnd), .vdd(vdd), .A(_12150_), .B(_12149_), .Y(_9805_) );
OAI21X1 OAI21X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_9798_), .B(_9802_), .C(_9805_), .Y(_9806_) );
NAND2X1 NAND2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_9804_), .B(_9806_), .Y(_9807_) );
NAND3X1 NAND3X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_9783_), .B(_9807_), .C(_9787_), .Y(_9808_) );
NAND3X1 NAND3X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_9351_), .B(_9774_), .C(_9778_), .Y(_9809_) );
NAND3X1 NAND3X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_9579_), .B(_9780_), .C(_9781_), .Y(_9810_) );
AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_9356_), .B(_9369_), .C(_9809_), .D(_9810_), .Y(_9811_) );
AOI21X1 AOI21X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_9779_), .B(_9782_), .C(_9578_), .Y(_9812_) );
INVX1 INVX1_1359 ( .gnd(gnd), .vdd(vdd), .A(_9807_), .Y(_9813_) );
OAI21X1 OAI21X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_9812_), .B(_9811_), .C(_9813_), .Y(_9814_) );
NAND3X1 NAND3X1_2197 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf2_), .B(_9814_), .C(_9808_), .Y(_9815_) );
INVX1 INVX1_1360 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf1_), .Y(_9816_) );
OAI21X1 OAI21X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_9812_), .B(_9811_), .C(_9807_), .Y(_9817_) );
NAND3X1 NAND3X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_9783_), .B(_9813_), .C(_9787_), .Y(_9818_) );
NAND3X1 NAND3X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_9816_), .B(_9817_), .C(_9818_), .Y(_9819_) );
NAND3X1 NAND3X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_9577_), .B(_9815_), .C(_9819_), .Y(_9820_) );
NAND3X1 NAND3X1_2201 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf0_), .B(_9817_), .C(_9818_), .Y(_9821_) );
NAND3X1 NAND3X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_9816_), .B(_9814_), .C(_9808_), .Y(_9822_) );
NAND3X1 NAND3X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_9372_), .B(_9821_), .C(_9822_), .Y(_9823_) );
NAND3X1 NAND3X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_9576_), .B(_9820_), .C(_9823_), .Y(_9824_) );
INVX1 INVX1_1361 ( .gnd(gnd), .vdd(vdd), .A(_9576_), .Y(_9825_) );
AOI21X1 AOI21X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_9821_), .B(_9822_), .C(_9372_), .Y(_9826_) );
AOI21X1 AOI21X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_9815_), .B(_9819_), .C(_9577_), .Y(_9827_) );
OAI21X1 OAI21X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_9826_), .B(_9827_), .C(_9825_), .Y(_9828_) );
INVX1 INVX1_1362 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf2_), .Y(_9829_) );
OAI21X1 OAI21X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_9798_), .B(_9802_), .C(_9829_), .Y(_9830_) );
NAND3X1 NAND3X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_9799_), .B(_9800_), .C(_9801_), .Y(_9831_) );
OAI21X1 OAI21X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_9794_), .B(_9797_), .C(_9131_), .Y(_9832_) );
NAND3X1 NAND3X1_2206 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf1_), .B(_9831_), .C(_9832_), .Y(_9833_) );
NAND2X1 NAND2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_9833_), .B(_9830_), .Y(_9834_) );
NOR2X1 NOR2X1_780 ( .gnd(gnd), .vdd(vdd), .A(_9134_), .B(_9834_), .Y(_9835_) );
INVX1 INVX1_1363 ( .gnd(gnd), .vdd(vdd), .A(_9134_), .Y(_9836_) );
AOI21X1 AOI21X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_9833_), .B(_9830_), .C(_9836_), .Y(_9837_) );
NOR3X1 NOR3X1_282 ( .gnd(gnd), .vdd(vdd), .A(_9137_), .B(_9837_), .C(_9835_), .Y(_9838_) );
NOR2X1 NOR2X1_781 ( .gnd(gnd), .vdd(vdd), .A(_8875_), .B(_9135_), .Y(_9839_) );
NAND3X1 NAND3X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_9830_), .B(_9833_), .C(_9836_), .Y(_9840_) );
INVX1 INVX1_1364 ( .gnd(gnd), .vdd(vdd), .A(_9837_), .Y(_9841_) );
AOI21X1 AOI21X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_9840_), .B(_9841_), .C(_9839_), .Y(_9842_) );
NOR2X1 NOR2X1_782 ( .gnd(gnd), .vdd(vdd), .A(_9842_), .B(_9838_), .Y(_9843_) );
OAI21X1 OAI21X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_12161_), .B(_12162_), .C(_9843_), .Y(_9844_) );
NOR2X1 NOR2X1_783 ( .gnd(gnd), .vdd(vdd), .A(_12162_), .B(_12161_), .Y(_9845_) );
OAI21X1 OAI21X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_9838_), .B(_9842_), .C(_9845_), .Y(_9846_) );
NAND2X1 NAND2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_9844_), .B(_9846_), .Y(_9847_) );
NAND3X1 NAND3X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9847_), .C(_9828_), .Y(_9848_) );
NAND3X1 NAND3X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_9372_), .B(_9815_), .C(_9819_), .Y(_9849_) );
NAND3X1 NAND3X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_9577_), .B(_9821_), .C(_9822_), .Y(_9850_) );
AOI21X1 AOI21X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_9849_), .B(_9850_), .C(_9825_), .Y(_9851_) );
AOI21X1 AOI21X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_9820_), .B(_9823_), .C(_9576_), .Y(_9852_) );
INVX1 INVX1_1365 ( .gnd(gnd), .vdd(vdd), .A(_9847_), .Y(_9853_) );
OAI21X1 OAI21X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_9851_), .B(_9852_), .C(_9853_), .Y(_9854_) );
NAND3X1 NAND3X1_2211 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_134_), .B(_9848_), .C(_9854_), .Y(_9855_) );
INVX1 INVX1_1366 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_134_), .Y(_9856_) );
NAND3X1 NAND3X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9853_), .C(_9828_), .Y(_9857_) );
OAI21X1 OAI21X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_9851_), .B(_9852_), .C(_9847_), .Y(_9858_) );
NAND3X1 NAND3X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_9856_), .B(_9857_), .C(_9858_), .Y(_9859_) );
NAND3X1 NAND3X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_9574_), .B(_9855_), .C(_9859_), .Y(_9860_) );
NAND3X1 NAND3X1_2215 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_134_), .B(_9857_), .C(_9858_), .Y(_9861_) );
NAND3X1 NAND3X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_9856_), .B(_9848_), .C(_9854_), .Y(_9862_) );
NAND3X1 NAND3X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_9399_), .B(_9861_), .C(_9862_), .Y(_9863_) );
NAND3X1 NAND3X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_9573_), .B(_9860_), .C(_9863_), .Y(_9864_) );
INVX2 INVX2_345 ( .gnd(gnd), .vdd(vdd), .A(_9573_), .Y(_9865_) );
AOI21X1 AOI21X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_9861_), .B(_9862_), .C(_9399_), .Y(_9866_) );
AOI21X1 AOI21X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_9855_), .B(_9859_), .C(_9574_), .Y(_9867_) );
OAI21X1 OAI21X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_9866_), .B(_9867_), .C(_9865_), .Y(_9868_) );
INVX1 INVX1_1367 ( .gnd(gnd), .vdd(vdd), .A(_9140_), .Y(_9869_) );
INVX1 INVX1_1368 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf0_), .Y(_9870_) );
OAI21X1 OAI21X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_9838_), .B(_9842_), .C(_9870_), .Y(_9871_) );
NAND3X1 NAND3X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_9839_), .B(_9840_), .C(_9841_), .Y(_9872_) );
OAI21X1 OAI21X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_9835_), .B(_9837_), .C(_9137_), .Y(_9873_) );
NAND3X1 NAND3X1_2220 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf4_), .B(_9873_), .C(_9872_), .Y(_9874_) );
NAND3X1 NAND3X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_9871_), .B(_9874_), .C(_9869_), .Y(_9875_) );
AOI21X1 AOI21X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_9873_), .B(_9872_), .C(bloque_datos_90_bF_buf3_), .Y(_9876_) );
NOR3X1 NOR3X1_283 ( .gnd(gnd), .vdd(vdd), .A(_9842_), .B(_9870_), .C(_9838_), .Y(_9877_) );
OAI21X1 OAI21X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_9877_), .B(_9876_), .C(_9140_), .Y(_9878_) );
AND2X2 AND2X2_217 ( .gnd(gnd), .vdd(vdd), .A(_9878_), .B(_9875_), .Y(_9879_) );
NAND2X1 NAND2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .B(_9879_), .Y(_9880_) );
INVX1 INVX1_1369 ( .gnd(gnd), .vdd(vdd), .A(_9880_), .Y(_9881_) );
NOR2X1 NOR2X1_784 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .B(_9879_), .Y(_9882_) );
NOR2X1 NOR2X1_785 ( .gnd(gnd), .vdd(vdd), .A(_9882_), .B(_9881_), .Y(_9883_) );
INVX4 INVX4_9 ( .gnd(gnd), .vdd(vdd), .A(_9883_), .Y(_9884_) );
NAND3X1 NAND3X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_9864_), .B(_9884_), .C(_9868_), .Y(_9885_) );
NAND3X1 NAND3X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_9399_), .B(_9855_), .C(_9859_), .Y(_9886_) );
NAND3X1 NAND3X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_9574_), .B(_9861_), .C(_9862_), .Y(_9887_) );
AOI21X1 AOI21X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_9886_), .B(_9887_), .C(_9865_), .Y(_9888_) );
AOI21X1 AOI21X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_9860_), .B(_9863_), .C(_9573_), .Y(_9889_) );
OAI21X1 OAI21X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_9888_), .B(_9889_), .C(_9883_), .Y(_9890_) );
NAND3X1 NAND3X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_9572_), .B(_9885_), .C(_9890_), .Y(_9891_) );
NAND2X1 NAND2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_150_), .B(_9891_), .Y(_9892_) );
INVX2 INVX2_346 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_150_), .Y(_9893_) );
OAI21X1 OAI21X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_9888_), .B(_9889_), .C(_9884_), .Y(_9894_) );
NAND3X1 NAND3X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_9864_), .B(_9883_), .C(_9868_), .Y(_9895_) );
AOI21X1 AOI21X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_9895_), .B(_9894_), .C(_9571_), .Y(_9896_) );
NAND2X1 NAND2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_9893_), .B(_9896_), .Y(_9897_) );
NAND3X1 NAND3X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_9422_), .B(_9892_), .C(_9897_), .Y(_9898_) );
NAND2X1 NAND2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_150_), .B(_9896_), .Y(_9899_) );
NAND2X1 NAND2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_9893_), .B(_9891_), .Y(_9900_) );
NAND3X1 NAND3X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_9416_), .B(_9900_), .C(_9899_), .Y(_9901_) );
AOI21X1 AOI21X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_9898_), .B(_9901_), .C(_9570_), .Y(_9902_) );
INVX1 INVX1_1370 ( .gnd(gnd), .vdd(vdd), .A(_9428_), .Y(_9903_) );
OAI21X1 OAI21X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_9903_), .B(_9220_), .C(_9427_), .Y(_9904_) );
NAND3X1 NAND3X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_9416_), .B(_9892_), .C(_9897_), .Y(_9905_) );
NAND3X1 NAND3X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_9422_), .B(_9900_), .C(_9899_), .Y(_9906_) );
AOI21X1 AOI21X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_9905_), .B(_9906_), .C(_9904_), .Y(_9907_) );
INVX1 INVX1_1371 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_138_), .Y(_9908_) );
OAI21X1 OAI21X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_9881_), .B(_9882_), .C(_9908_), .Y(_9909_) );
NAND2X1 NAND2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_138_), .B(_9883_), .Y(_9910_) );
NAND2X1 NAND2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_9909_), .B(_9910_), .Y(_9911_) );
NOR2X1 NOR2X1_786 ( .gnd(gnd), .vdd(vdd), .A(_9148_), .B(_9911_), .Y(_9912_) );
INVX1 INVX1_1372 ( .gnd(gnd), .vdd(vdd), .A(_9912_), .Y(_9913_) );
OAI21X1 OAI21X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_9086_), .B(_9145_), .C(_9911_), .Y(_9914_) );
NAND3X1 NAND3X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_9151_), .B(_9914_), .C(_9913_), .Y(_9915_) );
INVX1 INVX1_1373 ( .gnd(gnd), .vdd(vdd), .A(_9914_), .Y(_9916_) );
OAI21X1 OAI21X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_9916_), .B(_9912_), .C(_9152_), .Y(_9917_) );
NAND2X1 NAND2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_9917_), .B(_9915_), .Y(_9918_) );
INVX2 INVX2_347 ( .gnd(gnd), .vdd(vdd), .A(_9918_), .Y(_9919_) );
OAI21X1 OAI21X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_9902_), .B(_9907_), .C(_9919_), .Y(_9920_) );
NAND3X1 NAND3X1_2232 ( .gnd(gnd), .vdd(vdd), .A(_9905_), .B(_9906_), .C(_9904_), .Y(_9921_) );
AOI21X1 AOI21X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_9900_), .B(_9899_), .C(_9422_), .Y(_9922_) );
AOI21X1 AOI21X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_9892_), .B(_9897_), .C(_9416_), .Y(_9923_) );
OAI21X1 OAI21X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_9922_), .B(_9923_), .C(_9570_), .Y(_9924_) );
NAND3X1 NAND3X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_9918_), .B(_9921_), .C(_9924_), .Y(_9925_) );
NAND3X1 NAND3X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_12397_), .B(_9925_), .C(_9920_), .Y(_9926_) );
NAND2X1 NAND2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_166_), .B(_9926_), .Y(_9927_) );
INVX2 INVX2_348 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_166_), .Y(_9928_) );
NAND3X1 NAND3X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_9919_), .B(_9921_), .C(_9924_), .Y(_9929_) );
OAI21X1 OAI21X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_9902_), .B(_9907_), .C(_9918_), .Y(_9930_) );
AOI21X1 AOI21X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_9929_), .B(_9930_), .C(_12184_), .Y(_9931_) );
NAND2X1 NAND2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_9928_), .B(_9931_), .Y(_9932_) );
NAND3X1 NAND3X1_2236 ( .gnd(gnd), .vdd(vdd), .A(_9441_), .B(_9927_), .C(_9932_), .Y(_9933_) );
NAND2X1 NAND2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_166_), .B(_9931_), .Y(_9934_) );
NAND2X1 NAND2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_9928_), .B(_9926_), .Y(_9935_) );
NAND3X1 NAND3X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_9435_), .B(_9935_), .C(_9934_), .Y(_9936_) );
AOI21X1 AOI21X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_9933_), .B(_9936_), .C(_9568_), .Y(_9937_) );
NOR3X1 NOR3X1_284 ( .gnd(gnd), .vdd(vdd), .A(_9442_), .B(_9217_), .C(_9441_), .Y(_9938_) );
OAI21X1 OAI21X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_9938_), .B(_9216_), .C(_9446_), .Y(_9939_) );
NAND3X1 NAND3X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_9435_), .B(_9927_), .C(_9932_), .Y(_9940_) );
NAND3X1 NAND3X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_9441_), .B(_9935_), .C(_9934_), .Y(_9941_) );
AOI21X1 AOI21X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_9940_), .B(_9941_), .C(_9939_), .Y(_9942_) );
INVX1 INVX1_1374 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_154_), .Y(_9943_) );
NAND2X1 NAND2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_9943_), .B(_9918_), .Y(_9944_) );
NOR2X1 NOR2X1_787 ( .gnd(gnd), .vdd(vdd), .A(_9943_), .B(_9918_), .Y(_9945_) );
INVX2 INVX2_349 ( .gnd(gnd), .vdd(vdd), .A(_9945_), .Y(_9946_) );
NAND3X1 NAND3X1_2240 ( .gnd(gnd), .vdd(vdd), .A(_9155_), .B(_9944_), .C(_9946_), .Y(_9947_) );
INVX1 INVX1_1375 ( .gnd(gnd), .vdd(vdd), .A(_9944_), .Y(_9948_) );
OAI21X1 OAI21X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_9948_), .B(_9945_), .C(_9156_), .Y(_9949_) );
NAND3X1 NAND3X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_9159_), .B(_9949_), .C(_9947_), .Y(_9950_) );
NAND2X1 NAND2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_9949_), .B(_9947_), .Y(_9951_) );
OAI21X1 OAI21X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_9083_), .B(_9157_), .C(_9951_), .Y(_9952_) );
NAND2X1 NAND2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_9950_), .B(_9952_), .Y(_9953_) );
INVX1 INVX1_1376 ( .gnd(gnd), .vdd(vdd), .A(_9953_), .Y(_9954_) );
OAI21X1 OAI21X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_9937_), .B(_9942_), .C(_9954_), .Y(_9955_) );
NAND3X1 NAND3X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_9939_), .B(_9940_), .C(_9941_), .Y(_9956_) );
AOI21X1 AOI21X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_9935_), .B(_9934_), .C(_9441_), .Y(_9957_) );
AOI21X1 AOI21X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_9927_), .B(_9932_), .C(_9435_), .Y(_9958_) );
OAI21X1 OAI21X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_9957_), .B(_9958_), .C(_9568_), .Y(_9959_) );
NAND3X1 NAND3X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_9953_), .B(_9956_), .C(_9959_), .Y(_9960_) );
NAND3X1 NAND3X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_9566_), .B(_9960_), .C(_9955_), .Y(_9961_) );
NAND2X1 NAND2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_182_), .B(_9961_), .Y(_9962_) );
INVX2 INVX2_350 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_182_), .Y(_9963_) );
NAND3X1 NAND3X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_9954_), .B(_9956_), .C(_9959_), .Y(_9964_) );
OAI21X1 OAI21X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_9937_), .B(_9942_), .C(_9953_), .Y(_9965_) );
AOI21X1 AOI21X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_9964_), .B(_9965_), .C(_12194_), .Y(_9966_) );
NAND2X1 NAND2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_9963_), .B(_9966_), .Y(_9967_) );
NAND3X1 NAND3X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_9452_), .B(_9962_), .C(_9967_), .Y(_9968_) );
NAND2X1 NAND2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_9964_), .B(_9965_), .Y(_9969_) );
NAND3X1 NAND3X1_2247 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_182_), .B(_9566_), .C(_9969_), .Y(_9970_) );
NAND2X1 NAND2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_9963_), .B(_9961_), .Y(_9971_) );
NAND3X1 NAND3X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_9970_), .C(_9971_), .Y(_9972_) );
NAND3X1 NAND3X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_9972_), .B(_9565_), .C(_9968_), .Y(_9973_) );
AOI21X1 AOI21X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_9452_), .B(_9457_), .C(_8962_), .Y(_9974_) );
AOI21X1 AOI21X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_9465_), .B(_9463_), .C(_9974_), .Y(_9975_) );
AOI21X1 AOI21X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_9970_), .B(_9971_), .C(_9459_), .Y(_9976_) );
AOI21X1 AOI21X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_9962_), .B(_9967_), .C(_9452_), .Y(_9977_) );
OAI21X1 OAI21X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_9977_), .B(_9976_), .C(_9975_), .Y(_9978_) );
INVX1 INVX1_1377 ( .gnd(gnd), .vdd(vdd), .A(_9168_), .Y(_9979_) );
INVX1 INVX1_1378 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_170_), .Y(_9980_) );
NAND2X1 NAND2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_9980_), .B(_9953_), .Y(_9981_) );
INVX1 INVX1_1379 ( .gnd(gnd), .vdd(vdd), .A(_9981_), .Y(_9982_) );
NOR2X1 NOR2X1_788 ( .gnd(gnd), .vdd(vdd), .A(_9980_), .B(_9953_), .Y(_9983_) );
NOR2X1 NOR2X1_789 ( .gnd(gnd), .vdd(vdd), .A(_9983_), .B(_9982_), .Y(_9984_) );
AND2X2 AND2X2_218 ( .gnd(gnd), .vdd(vdd), .A(_9984_), .B(_9165_), .Y(_9985_) );
OAI21X1 OAI21X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_9982_), .B(_9983_), .C(_9164_), .Y(_9986_) );
INVX1 INVX1_1380 ( .gnd(gnd), .vdd(vdd), .A(_9986_), .Y(_9987_) );
NOR2X1 NOR2X1_790 ( .gnd(gnd), .vdd(vdd), .A(_9987_), .B(_9985_), .Y(_9988_) );
NAND2X1 NAND2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_9979_), .B(_9988_), .Y(_9989_) );
OAI21X1 OAI21X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_9985_), .B(_9987_), .C(_9168_), .Y(_9990_) );
NAND2X1 NAND2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_9990_), .B(_9989_), .Y(_9991_) );
NAND3X1 NAND3X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_9973_), .B(_9991_), .C(_9978_), .Y(_9992_) );
NAND3X1 NAND3X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_9962_), .C(_9967_), .Y(_9993_) );
NAND3X1 NAND3X1_2252 ( .gnd(gnd), .vdd(vdd), .A(_9452_), .B(_9970_), .C(_9971_), .Y(_9994_) );
AOI21X1 AOI21X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_9994_), .B(_9993_), .C(_9975_), .Y(_9995_) );
AOI21X1 AOI21X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_9972_), .B(_9968_), .C(_9565_), .Y(_9996_) );
INVX1 INVX1_1381 ( .gnd(gnd), .vdd(vdd), .A(_9991_), .Y(_9997_) );
OAI21X1 OAI21X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_9995_), .B(_9996_), .C(_9997_), .Y(_9998_) );
NAND3X1 NAND3X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_9563_), .B(_9992_), .C(_9998_), .Y(_9999_) );
NAND2X1 NAND2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_198_), .B(_9999_), .Y(_10000_) );
INVX2 INVX2_351 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_198_), .Y(_10001_) );
AOI21X1 AOI21X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_9973_), .B(_9978_), .C(_9991_), .Y(_10002_) );
NOR2X1 NOR2X1_791 ( .gnd(gnd), .vdd(vdd), .A(_9562_), .B(_10002_), .Y(_10003_) );
NAND3X1 NAND3X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_10001_), .B(_9992_), .C(_10003_), .Y(_10004_) );
NAND3X1 NAND3X1_2255 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_10000_), .C(_10004_), .Y(_10005_) );
NAND3X1 NAND3X1_2256 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_198_), .B(_9992_), .C(_10003_), .Y(_10006_) );
NAND2X1 NAND2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_10001_), .B(_9999_), .Y(_10007_) );
NAND3X1 NAND3X1_2257 ( .gnd(gnd), .vdd(vdd), .A(_9472_), .B(_10007_), .C(_10006_), .Y(_10008_) );
AOI21X1 AOI21X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_10005_), .B(_10008_), .C(_9561_), .Y(_10009_) );
NOR3X1 NOR3X1_285 ( .gnd(gnd), .vdd(vdd), .A(_9479_), .B(_9211_), .C(_9478_), .Y(_10010_) );
OAI21X1 OAI21X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_10010_), .B(_9210_), .C(_9483_), .Y(_10011_) );
NAND3X1 NAND3X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_9472_), .B(_10000_), .C(_10004_), .Y(_10012_) );
NAND3X1 NAND3X1_2259 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_10007_), .C(_10006_), .Y(_10013_) );
AOI21X1 AOI21X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_10012_), .B(_10013_), .C(_10011_), .Y(_10014_) );
INVX1 INVX1_1382 ( .gnd(gnd), .vdd(vdd), .A(_9176_), .Y(_10015_) );
INVX1 INVX1_1383 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_186_), .Y(_10016_) );
NAND2X1 NAND2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_10016_), .B(_9991_), .Y(_10017_) );
NOR2X1 NOR2X1_792 ( .gnd(gnd), .vdd(vdd), .A(_10016_), .B(_9991_), .Y(_10018_) );
INVX1 INVX1_1384 ( .gnd(gnd), .vdd(vdd), .A(_10018_), .Y(_10019_) );
NAND3X1 NAND3X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_9173_), .B(_10017_), .C(_10019_), .Y(_10020_) );
INVX1 INVX1_1385 ( .gnd(gnd), .vdd(vdd), .A(_10017_), .Y(_10021_) );
OAI21X1 OAI21X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_10021_), .B(_10018_), .C(_9172_), .Y(_10022_) );
NAND3X1 NAND3X1_2261 ( .gnd(gnd), .vdd(vdd), .A(_10015_), .B(_10022_), .C(_10020_), .Y(_10023_) );
INVX1 INVX1_1386 ( .gnd(gnd), .vdd(vdd), .A(_10020_), .Y(_10024_) );
INVX1 INVX1_1387 ( .gnd(gnd), .vdd(vdd), .A(_10022_), .Y(_10025_) );
OAI21X1 OAI21X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_10024_), .B(_10025_), .C(_9176_), .Y(_10026_) );
NAND2X1 NAND2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_10023_), .B(_10026_), .Y(_10027_) );
INVX1 INVX1_1388 ( .gnd(gnd), .vdd(vdd), .A(_10027_), .Y(_10028_) );
OAI21X1 OAI21X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_10009_), .B(_10014_), .C(_10028_), .Y(_10029_) );
NAND3X1 NAND3X1_2262 ( .gnd(gnd), .vdd(vdd), .A(_10012_), .B(_10013_), .C(_10011_), .Y(_10030_) );
AOI21X1 AOI21X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_10007_), .B(_10006_), .C(_9478_), .Y(_10031_) );
AOI21X1 AOI21X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_10000_), .B(_10004_), .C(_9472_), .Y(_10032_) );
OAI21X1 OAI21X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_10031_), .B(_10032_), .C(_9561_), .Y(_10033_) );
NAND3X1 NAND3X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_10030_), .B(_10027_), .C(_10033_), .Y(_10034_) );
NAND3X1 NAND3X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_9559_), .B(_10034_), .C(_10029_), .Y(_10035_) );
NAND2X1 NAND2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_214_), .B(_10035_), .Y(_10036_) );
INVX2 INVX2_352 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_214_), .Y(_10037_) );
OAI21X1 OAI21X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_10009_), .B(_10014_), .C(_10027_), .Y(_10038_) );
NAND3X1 NAND3X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_10030_), .B(_10028_), .C(_10033_), .Y(_10039_) );
AOI21X1 AOI21X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_10039_), .B(_10038_), .C(_12212_), .Y(_10040_) );
NAND2X1 NAND2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_10037_), .B(_10040_), .Y(_10041_) );
NAND3X1 NAND3X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_9497_), .B(_10036_), .C(_10041_), .Y(_10042_) );
NAND2X1 NAND2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_214_), .B(_10040_), .Y(_10043_) );
NAND2X1 NAND2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_10037_), .B(_10035_), .Y(_10044_) );
NAND3X1 NAND3X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_9491_), .B(_10044_), .C(_10043_), .Y(_10045_) );
AOI21X1 AOI21X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_10042_), .B(_10045_), .C(_9558_), .Y(_10046_) );
NOR3X1 NOR3X1_286 ( .gnd(gnd), .vdd(vdd), .A(_9498_), .B(_9208_), .C(_9497_), .Y(_10047_) );
OAI21X1 OAI21X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_10047_), .B(_9207_), .C(_9502_), .Y(_10048_) );
NAND3X1 NAND3X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_9491_), .B(_10036_), .C(_10041_), .Y(_10049_) );
NAND3X1 NAND3X1_2269 ( .gnd(gnd), .vdd(vdd), .A(_9497_), .B(_10044_), .C(_10043_), .Y(_10050_) );
AOI21X1 AOI21X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_10049_), .B(_10050_), .C(_10048_), .Y(_10051_) );
INVX1 INVX1_1389 ( .gnd(gnd), .vdd(vdd), .A(_9184_), .Y(_10052_) );
INVX1 INVX1_1390 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_202_), .Y(_10053_) );
NAND2X1 NAND2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_10053_), .B(_10027_), .Y(_10054_) );
NOR2X1 NOR2X1_793 ( .gnd(gnd), .vdd(vdd), .A(_10053_), .B(_10027_), .Y(_10055_) );
INVX2 INVX2_353 ( .gnd(gnd), .vdd(vdd), .A(_10055_), .Y(_10056_) );
NAND3X1 NAND3X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_9181_), .B(_10054_), .C(_10056_), .Y(_10057_) );
INVX1 INVX1_1391 ( .gnd(gnd), .vdd(vdd), .A(_10054_), .Y(_10058_) );
OAI21X1 OAI21X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_10058_), .B(_10055_), .C(_9180_), .Y(_10059_) );
NAND3X1 NAND3X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_10052_), .B(_10059_), .C(_10057_), .Y(_10060_) );
INVX1 INVX1_1392 ( .gnd(gnd), .vdd(vdd), .A(_10057_), .Y(_10061_) );
INVX1 INVX1_1393 ( .gnd(gnd), .vdd(vdd), .A(_10059_), .Y(_10062_) );
OAI21X1 OAI21X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_10061_), .B(_10062_), .C(_9184_), .Y(_10063_) );
NAND2X1 NAND2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_10060_), .B(_10063_), .Y(_10064_) );
INVX2 INVX2_354 ( .gnd(gnd), .vdd(vdd), .A(_10064_), .Y(_10065_) );
OAI21X1 OAI21X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_10051_), .B(_10046_), .C(_10065_), .Y(_10066_) );
NAND3X1 NAND3X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_10049_), .B(_10050_), .C(_10048_), .Y(_10067_) );
AOI21X1 AOI21X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_10044_), .B(_10043_), .C(_9497_), .Y(_10068_) );
AOI21X1 AOI21X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10041_), .C(_9491_), .Y(_10069_) );
OAI21X1 OAI21X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_10068_), .B(_10069_), .C(_9558_), .Y(_10070_) );
NAND3X1 NAND3X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_10064_), .B(_10070_), .C(_10067_), .Y(_10071_) );
NAND3X1 NAND3X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_9556_), .B(_10071_), .C(_10066_), .Y(_10072_) );
NAND2X1 NAND2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_230_), .B(_10072_), .Y(_10073_) );
INVX2 INVX2_355 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_230_), .Y(_10074_) );
OAI21X1 OAI21X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_10051_), .B(_10046_), .C(_10064_), .Y(_10075_) );
NAND3X1 NAND3X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_10065_), .B(_10070_), .C(_10067_), .Y(_10076_) );
AOI21X1 AOI21X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_10076_), .B(_10075_), .C(_9555_), .Y(_10077_) );
NAND2X1 NAND2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_10074_), .B(_10077_), .Y(_10078_) );
NAND3X1 NAND3X1_2276 ( .gnd(gnd), .vdd(vdd), .A(_9516_), .B(_10073_), .C(_10078_), .Y(_10079_) );
NAND2X1 NAND2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_230_), .B(_10077_), .Y(_10080_) );
NAND2X1 NAND2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_10074_), .B(_10072_), .Y(_10081_) );
NAND3X1 NAND3X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_9510_), .B(_10081_), .C(_10080_), .Y(_10082_) );
AOI21X1 AOI21X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_10079_), .B(_10082_), .C(_9552_), .Y(_10083_) );
NOR3X1 NOR3X1_287 ( .gnd(gnd), .vdd(vdd), .A(_9517_), .B(_9205_), .C(_9516_), .Y(_10084_) );
OAI21X1 OAI21X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_10084_), .B(_9204_), .C(_9521_), .Y(_10085_) );
NAND3X1 NAND3X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_9510_), .B(_10073_), .C(_10078_), .Y(_10086_) );
NAND3X1 NAND3X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_9516_), .B(_10081_), .C(_10080_), .Y(_10087_) );
AOI21X1 AOI21X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_10086_), .B(_10087_), .C(_10085_), .Y(_10088_) );
INVX1 INVX1_1394 ( .gnd(gnd), .vdd(vdd), .A(_9192_), .Y(_10089_) );
INVX1 INVX1_1395 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_218_), .Y(_10090_) );
NAND2X1 NAND2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_10090_), .B(_10064_), .Y(_10091_) );
NOR2X1 NOR2X1_794 ( .gnd(gnd), .vdd(vdd), .A(_10090_), .B(_10064_), .Y(_10092_) );
INVX2 INVX2_356 ( .gnd(gnd), .vdd(vdd), .A(_10092_), .Y(_10093_) );
NAND2X1 NAND2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_10091_), .B(_10093_), .Y(_10094_) );
OR2X2 OR2X2_236 ( .gnd(gnd), .vdd(vdd), .A(_10094_), .B(_9188_), .Y(_10095_) );
AOI21X1 AOI21X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_10091_), .B(_10093_), .C(_9189_), .Y(_10096_) );
INVX1 INVX1_1396 ( .gnd(gnd), .vdd(vdd), .A(_10096_), .Y(_10097_) );
NAND3X1 NAND3X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_10089_), .B(_10097_), .C(_10095_), .Y(_10098_) );
NOR2X1 NOR2X1_795 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .B(_10094_), .Y(_10099_) );
OAI21X1 OAI21X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_10099_), .B(_10096_), .C(_9192_), .Y(_10100_) );
NAND2X1 NAND2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_10100_), .B(_10098_), .Y(_10101_) );
INVX2 INVX2_357 ( .gnd(gnd), .vdd(vdd), .A(_10101_), .Y(_10102_) );
OAI21X1 OAI21X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_10088_), .B(_10083_), .C(_10102_), .Y(_10103_) );
NAND3X1 NAND3X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_10086_), .B(_10087_), .C(_10085_), .Y(_10104_) );
AOI21X1 AOI21X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_10081_), .B(_10080_), .C(_9516_), .Y(_10105_) );
AOI21X1 AOI21X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_10073_), .B(_10078_), .C(_9510_), .Y(_10106_) );
OAI21X1 OAI21X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_10105_), .B(_10106_), .C(_9552_), .Y(_10107_) );
NAND3X1 NAND3X1_2282 ( .gnd(gnd), .vdd(vdd), .A(_10107_), .B(_10101_), .C(_10104_), .Y(_10108_) );
NAND3X1 NAND3X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_12462_), .B(_10108_), .C(_10103_), .Y(_10109_) );
NAND2X1 NAND2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_246_), .B(_10109_), .Y(_10110_) );
INVX1 INVX1_1397 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_246_), .Y(_10111_) );
NAND3X1 NAND3X1_2284 ( .gnd(gnd), .vdd(vdd), .A(_10107_), .B(_10102_), .C(_10104_), .Y(_10112_) );
OAI21X1 OAI21X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_10088_), .B(_10083_), .C(_10101_), .Y(_10113_) );
AOI21X1 AOI21X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_10112_), .B(_10113_), .C(_12234_), .Y(_10114_) );
NAND2X1 NAND2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_10111_), .B(_10114_), .Y(_10115_) );
NAND3X1 NAND3X1_2285 ( .gnd(gnd), .vdd(vdd), .A(_9535_), .B(_10110_), .C(_10115_), .Y(_10116_) );
NAND2X1 NAND2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_246_), .B(_10114_), .Y(_10117_) );
NAND2X1 NAND2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_10111_), .B(_10109_), .Y(_10118_) );
NAND3X1 NAND3X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_9527_), .B(_10118_), .C(_10117_), .Y(_10119_) );
AOI21X1 AOI21X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_10116_), .B(_10119_), .C(_9550_), .Y(_10120_) );
OAI21X1 OAI21X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_9540_), .B(_9539_), .C(_9537_), .Y(_10121_) );
NAND3X1 NAND3X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_9527_), .B(_10110_), .C(_10115_), .Y(_10122_) );
NAND3X1 NAND3X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_9535_), .B(_10118_), .C(_10117_), .Y(_10123_) );
AOI21X1 AOI21X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_10122_), .B(_10123_), .C(_10121_), .Y(_10124_) );
INVX1 INVX1_1398 ( .gnd(gnd), .vdd(vdd), .A(_9200_), .Y(_10125_) );
NOR2X1 NOR2X1_796 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_234_), .B(_10102_), .Y(_10126_) );
INVX1 INVX1_1399 ( .gnd(gnd), .vdd(vdd), .A(_10126_), .Y(_10127_) );
NAND2X1 NAND2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_234_), .B(_10102_), .Y(_10128_) );
NAND3X1 NAND3X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_10128_), .C(_10127_), .Y(_10129_) );
INVX2 INVX2_358 ( .gnd(gnd), .vdd(vdd), .A(_10128_), .Y(_10130_) );
OAI21X1 OAI21X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_10130_), .B(_10126_), .C(_9196_), .Y(_10131_) );
NAND3X1 NAND3X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_10125_), .B(_10131_), .C(_10129_), .Y(_10132_) );
NOR3X1 NOR3X1_288 ( .gnd(gnd), .vdd(vdd), .A(_9196_), .B(_10126_), .C(_10130_), .Y(_10133_) );
AOI21X1 AOI21X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_10128_), .B(_10127_), .C(_9197_), .Y(_10134_) );
OAI21X1 OAI21X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_10134_), .B(_10133_), .C(_9200_), .Y(_10135_) );
NAND2X1 NAND2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_10132_), .B(_10135_), .Y(_10136_) );
INVX2 INVX2_359 ( .gnd(gnd), .vdd(vdd), .A(_10136_), .Y(_10137_) );
OAI21X1 OAI21X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_10124_), .B(_10120_), .C(_10137_), .Y(_10138_) );
NAND3X1 NAND3X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_10122_), .B(_10123_), .C(_10121_), .Y(_10139_) );
NAND3X1 NAND3X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_10116_), .B(_10119_), .C(_9550_), .Y(_10140_) );
NAND3X1 NAND3X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_10140_), .B(_10136_), .C(_10139_), .Y(_10141_) );
NAND2X1 NAND2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_10141_), .B(_10138_), .Y(_10142_) );
XOR2X1 XOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_10142_), .B(_9549_), .Y(module_2_H_6_) );
OAI21X1 OAI21X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_10124_), .B(_10120_), .C(_10136_), .Y(_10143_) );
NAND3X1 NAND3X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_10140_), .B(_10137_), .C(_10139_), .Y(_10144_) );
NAND3X1 NAND3X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_10144_), .B(_10143_), .C(_9549_), .Y(_10145_) );
AOI21X1 AOI21X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_10118_), .B(_10117_), .C(_9535_), .Y(_10146_) );
AOI21X1 AOI21X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_10123_), .B(_10121_), .C(_10146_), .Y(_10147_) );
AOI21X1 AOI21X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_10125_), .B(_10131_), .C(_10133_), .Y(_10148_) );
OAI21X1 OAI21X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_9192_), .B(_10096_), .C(_10095_), .Y(_10149_) );
AOI21X1 AOI21X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_10052_), .B(_10059_), .C(_10061_), .Y(_10150_) );
INVX1 INVX1_1400 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_203_), .Y(_10151_) );
OAI21X1 OAI21X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_10025_), .B(_9176_), .C(_10020_), .Y(_10152_) );
INVX1 INVX1_1401 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_187_), .Y(_10153_) );
AOI21X1 AOI21X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_9979_), .B(_9986_), .C(_9985_), .Y(_10154_) );
INVX1 INVX1_1402 ( .gnd(gnd), .vdd(vdd), .A(_10154_), .Y(_10155_) );
INVX1 INVX1_1403 ( .gnd(gnd), .vdd(vdd), .A(_9983_), .Y(_10156_) );
INVX1 INVX1_1404 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_171_), .Y(_10157_) );
OAI21X1 OAI21X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_9951_), .B(_9160_), .C(_9947_), .Y(_10158_) );
INVX1 INVX1_1405 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_155_), .Y(_10159_) );
AOI21X1 AOI21X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_9151_), .B(_9914_), .C(_9912_), .Y(_10160_) );
INVX1 INVX1_1406 ( .gnd(gnd), .vdd(vdd), .A(_9878_), .Y(_10161_) );
OAI21X1 OAI21X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_10161_), .B(_9144_), .C(_9875_), .Y(_10162_) );
OAI21X1 OAI21X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_9137_), .B(_9837_), .C(_9840_), .Y(_10163_) );
INVX1 INVX1_1407 ( .gnd(gnd), .vdd(vdd), .A(_9833_), .Y(_10164_) );
OAI21X1 OAI21X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_9131_), .B(_9797_), .C(_9800_), .Y(_10165_) );
AOI21X1 AOI21X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_9758_), .B(_9760_), .C(_9753_), .Y(_10166_) );
INVX1 INVX1_1408 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf1_), .Y(_10167_) );
NOR2X1 NOR2X1_797 ( .gnd(gnd), .vdd(vdd), .A(_9093_), .B(_9114_), .Y(_10168_) );
AOI21X1 AOI21X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_10168_), .B(_9717_), .C(_9720_), .Y(_10169_) );
INVX1 INVX1_1409 ( .gnd(gnd), .vdd(vdd), .A(_9681_), .Y(_10170_) );
AOI21X1 AOI21X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_9674_), .B(_10170_), .C(_9680_), .Y(_10171_) );
INVX1 INVX1_1410 ( .gnd(gnd), .vdd(vdd), .A(_9678_), .Y(_10172_) );
INVX1 INVX1_1411 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .Y(_10173_) );
OAI21X1 OAI21X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_9648_), .B(_9645_), .C(_9641_), .Y(_10174_) );
NOR2X1 NOR2X1_798 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_27_), .B(module_2_W_11_), .Y(_10175_) );
INVX1 INVX1_1412 ( .gnd(gnd), .vdd(vdd), .A(_10175_), .Y(_10176_) );
NAND2X1 NAND2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_27_), .B(module_2_W_11_), .Y(_10177_) );
NAND2X1 NAND2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_10177_), .B(_10176_), .Y(_10178_) );
NAND3X1 NAND3X1_2296 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_26_), .B(module_2_W_10_), .C(_10178_), .Y(_10179_) );
NAND3X1 NAND3X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_9637_), .B(_10177_), .C(_10176_), .Y(_10180_) );
NAND2X1 NAND2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_10180_), .B(_10179_), .Y(_10181_) );
XOR2X1 XOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_10174_), .B(_10181_), .Y(_10182_) );
NAND2X1 NAND2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_10173_), .B(_10182_), .Y(_10183_) );
XNOR2X1 XNOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_10174_), .B(_10181_), .Y(_10184_) );
NAND2X1 NAND2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .B(_10184_), .Y(_10185_) );
NAND2X1 NAND2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_10185_), .B(_10183_), .Y(_10186_) );
NAND2X1 NAND2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_10172_), .B(_10186_), .Y(_10187_) );
NAND3X1 NAND3X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_9678_), .B(_10185_), .C(_10183_), .Y(_10188_) );
NAND2X1 NAND2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_10188_), .B(_10187_), .Y(_10189_) );
XNOR2X1 XNOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_10189_), .B(_10171_), .Y(_10190_) );
NAND2X1 NAND2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf0_), .B(_10190_), .Y(_10191_) );
INVX1 INVX1_1413 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf4_), .Y(_10192_) );
OR2X2 OR2X2_237 ( .gnd(gnd), .vdd(vdd), .A(_9679_), .B(_9675_), .Y(_10193_) );
OAI21X1 OAI21X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_9109_), .B(_9681_), .C(_10193_), .Y(_10194_) );
XNOR2X1 XNOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_10189_), .B(_10194_), .Y(_10195_) );
NAND2X1 NAND2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_10192_), .B(_10195_), .Y(_10196_) );
NAND2X1 NAND2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_10191_), .B(_10196_), .Y(_10197_) );
NOR2X1 NOR2X1_799 ( .gnd(gnd), .vdd(vdd), .A(_9712_), .B(_10197_), .Y(_10198_) );
AOI21X1 AOI21X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_10191_), .B(_10196_), .C(_9716_), .Y(_10199_) );
OAI21X1 OAI21X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_10198_), .B(_10199_), .C(_10169_), .Y(_10200_) );
OAI21X1 OAI21X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_9721_), .B(_9115_), .C(_9713_), .Y(_10201_) );
OR2X2 OR2X2_238 ( .gnd(gnd), .vdd(vdd), .A(_10197_), .B(_9712_), .Y(_10202_) );
INVX1 INVX1_1414 ( .gnd(gnd), .vdd(vdd), .A(_10199_), .Y(_10203_) );
NAND3X1 NAND3X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_10203_), .B(_10201_), .C(_10202_), .Y(_10204_) );
NAND2X1 NAND2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_10200_), .B(_10204_), .Y(_10205_) );
NAND2X1 NAND2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_10167_), .B(_10205_), .Y(_10206_) );
AND2X2 AND2X2_219 ( .gnd(gnd), .vdd(vdd), .A(_10204_), .B(_10200_), .Y(_10207_) );
NAND2X1 NAND2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf0_), .B(_10207_), .Y(_10208_) );
AOI21X1 AOI21X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_10206_), .B(_10208_), .C(_9755_), .Y(_10209_) );
NAND3X1 NAND3X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_9755_), .B(_10206_), .C(_10208_), .Y(_10210_) );
INVX2 INVX2_360 ( .gnd(gnd), .vdd(vdd), .A(_10210_), .Y(_10211_) );
OAI21X1 OAI21X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_10211_), .B(_10209_), .C(_10166_), .Y(_10212_) );
INVX2 INVX2_361 ( .gnd(gnd), .vdd(vdd), .A(_10212_), .Y(_10213_) );
NOR2X1 NOR2X1_800 ( .gnd(gnd), .vdd(vdd), .A(_10209_), .B(_10211_), .Y(_10214_) );
OAI21X1 OAI21X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_9753_), .B(_9757_), .C(_10214_), .Y(_10215_) );
INVX2 INVX2_362 ( .gnd(gnd), .vdd(vdd), .A(_10215_), .Y(_10216_) );
OAI21X1 OAI21X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_10216_), .B(_10213_), .C(bloque_datos_59_bF_buf2_), .Y(_10217_) );
INVX1 INVX1_1415 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf1_), .Y(_10218_) );
NAND3X1 NAND3X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_10218_), .B(_10212_), .C(_10215_), .Y(_10219_) );
NAND3X1 NAND3X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_9793_), .B(_10219_), .C(_10217_), .Y(_10220_) );
OAI21X1 OAI21X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_10216_), .B(_10213_), .C(_10218_), .Y(_10221_) );
NAND3X1 NAND3X1_2303 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf0_), .B(_10212_), .C(_10215_), .Y(_10222_) );
NAND3X1 NAND3X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_9796_), .B(_10222_), .C(_10221_), .Y(_10223_) );
AOI21X1 AOI21X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_10220_), .B(_10223_), .C(_10165_), .Y(_10224_) );
NAND3X1 NAND3X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_10165_), .B(_10220_), .C(_10223_), .Y(_10225_) );
INVX2 INVX2_363 ( .gnd(gnd), .vdd(vdd), .A(_10225_), .Y(_10226_) );
OAI21X1 OAI21X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_10226_), .B(_10224_), .C(bloque_datos_75_bF_buf0_), .Y(_10227_) );
INVX1 INVX1_1416 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf4_), .Y(_10228_) );
INVX1 INVX1_1417 ( .gnd(gnd), .vdd(vdd), .A(_10224_), .Y(_10229_) );
NAND3X1 NAND3X1_2306 ( .gnd(gnd), .vdd(vdd), .A(_10228_), .B(_10225_), .C(_10229_), .Y(_10230_) );
NAND3X1 NAND3X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_10164_), .B(_10230_), .C(_10227_), .Y(_10231_) );
OAI21X1 OAI21X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_10226_), .B(_10224_), .C(_10228_), .Y(_10232_) );
NAND3X1 NAND3X1_2308 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf3_), .B(_10225_), .C(_10229_), .Y(_10233_) );
NAND3X1 NAND3X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_9833_), .B(_10233_), .C(_10232_), .Y(_10234_) );
AOI21X1 AOI21X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_10231_), .B(_10234_), .C(_10163_), .Y(_10235_) );
NAND3X1 NAND3X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_10163_), .B(_10231_), .C(_10234_), .Y(_10236_) );
INVX2 INVX2_364 ( .gnd(gnd), .vdd(vdd), .A(_10236_), .Y(_10237_) );
OAI21X1 OAI21X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_10237_), .B(_10235_), .C(bloque_datos_91_bF_buf1_), .Y(_10238_) );
INVX1 INVX1_1418 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf0_), .Y(_10239_) );
INVX1 INVX1_1419 ( .gnd(gnd), .vdd(vdd), .A(_10235_), .Y(_10240_) );
NAND3X1 NAND3X1_2311 ( .gnd(gnd), .vdd(vdd), .A(_10239_), .B(_10236_), .C(_10240_), .Y(_10241_) );
NAND3X1 NAND3X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_9877_), .B(_10241_), .C(_10238_), .Y(_10242_) );
OAI21X1 OAI21X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_10237_), .B(_10235_), .C(_10239_), .Y(_10243_) );
NAND3X1 NAND3X1_2313 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf3_), .B(_10236_), .C(_10240_), .Y(_10244_) );
NAND3X1 NAND3X1_2314 ( .gnd(gnd), .vdd(vdd), .A(_9874_), .B(_10244_), .C(_10243_), .Y(_10245_) );
NAND3X1 NAND3X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_10242_), .B(_10245_), .C(_10162_), .Y(_10246_) );
INVX1 INVX1_1420 ( .gnd(gnd), .vdd(vdd), .A(_10246_), .Y(_10247_) );
AOI21X1 AOI21X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_10242_), .B(_10245_), .C(_10162_), .Y(_10248_) );
NOR2X1 NOR2X1_801 ( .gnd(gnd), .vdd(vdd), .A(_10248_), .B(_10247_), .Y(_10249_) );
XNOR2X1 XNOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_10249_), .B(module_2_W_139_), .Y(_10250_) );
NOR2X1 NOR2X1_802 ( .gnd(gnd), .vdd(vdd), .A(_9910_), .B(_10250_), .Y(_10251_) );
INVX1 INVX1_1421 ( .gnd(gnd), .vdd(vdd), .A(_10251_), .Y(_10252_) );
OAI21X1 OAI21X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_9908_), .B(_9884_), .C(_10250_), .Y(_10253_) );
NAND2X1 NAND2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_10253_), .B(_10252_), .Y(_10254_) );
OR2X2 OR2X2_239 ( .gnd(gnd), .vdd(vdd), .A(_10254_), .B(_10160_), .Y(_10255_) );
INVX1 INVX1_1422 ( .gnd(gnd), .vdd(vdd), .A(_10253_), .Y(_10256_) );
OAI21X1 OAI21X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_10256_), .B(_10251_), .C(_10160_), .Y(_10257_) );
NAND2X1 NAND2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_10257_), .B(_10255_), .Y(_10258_) );
NAND2X1 NAND2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_10159_), .B(_10258_), .Y(_10259_) );
INVX1 INVX1_1423 ( .gnd(gnd), .vdd(vdd), .A(_10259_), .Y(_10260_) );
NOR2X1 NOR2X1_803 ( .gnd(gnd), .vdd(vdd), .A(_10159_), .B(_10258_), .Y(_10261_) );
NOR3X1 NOR3X1_289 ( .gnd(gnd), .vdd(vdd), .A(_9946_), .B(_10261_), .C(_10260_), .Y(_10262_) );
INVX2 INVX2_365 ( .gnd(gnd), .vdd(vdd), .A(_10261_), .Y(_10263_) );
AOI21X1 AOI21X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_10259_), .B(_10263_), .C(_9945_), .Y(_10264_) );
NOR2X1 NOR2X1_804 ( .gnd(gnd), .vdd(vdd), .A(_10262_), .B(_10264_), .Y(_10265_) );
AND2X2 AND2X2_220 ( .gnd(gnd), .vdd(vdd), .A(_10265_), .B(_10158_), .Y(_10266_) );
AND2X2 AND2X2_221 ( .gnd(gnd), .vdd(vdd), .A(_9950_), .B(_9947_), .Y(_10267_) );
OAI21X1 OAI21X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_10264_), .B(_10262_), .C(_10267_), .Y(_10268_) );
INVX2 INVX2_366 ( .gnd(gnd), .vdd(vdd), .A(_10268_), .Y(_10269_) );
OAI21X1 OAI21X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_10266_), .B(_10269_), .C(_10157_), .Y(_10270_) );
NOR2X1 NOR2X1_805 ( .gnd(gnd), .vdd(vdd), .A(_10269_), .B(_10266_), .Y(_10271_) );
NAND2X1 NAND2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_171_), .B(_10271_), .Y(_10272_) );
NAND2X1 NAND2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_10270_), .B(_10272_), .Y(_10273_) );
NOR2X1 NOR2X1_806 ( .gnd(gnd), .vdd(vdd), .A(_10156_), .B(_10273_), .Y(_10274_) );
AOI21X1 AOI21X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_10270_), .B(_10272_), .C(_9983_), .Y(_10275_) );
NOR2X1 NOR2X1_807 ( .gnd(gnd), .vdd(vdd), .A(_10275_), .B(_10274_), .Y(_10276_) );
AND2X2 AND2X2_222 ( .gnd(gnd), .vdd(vdd), .A(_10276_), .B(_10155_), .Y(_10277_) );
OAI21X1 OAI21X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_10274_), .B(_10275_), .C(_10154_), .Y(_10278_) );
INVX2 INVX2_367 ( .gnd(gnd), .vdd(vdd), .A(_10278_), .Y(_10279_) );
OAI21X1 OAI21X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_10277_), .B(_10279_), .C(_10153_), .Y(_10280_) );
NOR2X1 NOR2X1_808 ( .gnd(gnd), .vdd(vdd), .A(_10279_), .B(_10277_), .Y(_10281_) );
NAND2X1 NAND2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_187_), .B(_10281_), .Y(_10282_) );
NAND3X1 NAND3X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_10018_), .B(_10280_), .C(_10282_), .Y(_10283_) );
INVX2 INVX2_368 ( .gnd(gnd), .vdd(vdd), .A(_10283_), .Y(_10284_) );
AOI21X1 AOI21X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_10280_), .B(_10282_), .C(_10018_), .Y(_10285_) );
NOR2X1 NOR2X1_809 ( .gnd(gnd), .vdd(vdd), .A(_10285_), .B(_10284_), .Y(_10286_) );
NAND2X1 NAND2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_10152_), .B(_10286_), .Y(_10287_) );
AOI21X1 AOI21X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_10015_), .B(_10022_), .C(_10024_), .Y(_10288_) );
OAI21X1 OAI21X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_10284_), .B(_10285_), .C(_10288_), .Y(_10289_) );
NAND2X1 NAND2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_10289_), .B(_10287_), .Y(_10290_) );
NAND2X1 NAND2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_10151_), .B(_10290_), .Y(_10291_) );
NOR2X1 NOR2X1_810 ( .gnd(gnd), .vdd(vdd), .A(_10151_), .B(_10290_), .Y(_10292_) );
INVX2 INVX2_369 ( .gnd(gnd), .vdd(vdd), .A(_10292_), .Y(_10293_) );
NAND3X1 NAND3X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_10055_), .B(_10291_), .C(_10293_), .Y(_10294_) );
INVX1 INVX1_1424 ( .gnd(gnd), .vdd(vdd), .A(_10291_), .Y(_10295_) );
OAI21X1 OAI21X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_10295_), .B(_10292_), .C(_10056_), .Y(_10296_) );
NAND2X1 NAND2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_10296_), .B(_10294_), .Y(_10297_) );
NOR2X1 NOR2X1_811 ( .gnd(gnd), .vdd(vdd), .A(_10150_), .B(_10297_), .Y(_10298_) );
OAI21X1 OAI21X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_10062_), .B(_9184_), .C(_10057_), .Y(_10299_) );
AOI21X1 AOI21X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_10296_), .B(_10294_), .C(_10299_), .Y(_10300_) );
NOR2X1 NOR2X1_812 ( .gnd(gnd), .vdd(vdd), .A(_10300_), .B(_10298_), .Y(_10301_) );
NOR2X1 NOR2X1_813 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_219_), .B(_10301_), .Y(_10302_) );
AND2X2 AND2X2_223 ( .gnd(gnd), .vdd(vdd), .A(_10301_), .B(module_2_W_219_), .Y(_10303_) );
NOR3X1 NOR3X1_290 ( .gnd(gnd), .vdd(vdd), .A(_10302_), .B(_10093_), .C(_10303_), .Y(_10304_) );
OR2X2 OR2X2_240 ( .gnd(gnd), .vdd(vdd), .A(_10301_), .B(module_2_W_219_), .Y(_10305_) );
NAND2X1 NAND2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_219_), .B(_10301_), .Y(_10306_) );
AOI21X1 AOI21X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_10306_), .B(_10305_), .C(_10092_), .Y(_10307_) );
NOR2X1 NOR2X1_814 ( .gnd(gnd), .vdd(vdd), .A(_10307_), .B(_10304_), .Y(_10308_) );
AND2X2 AND2X2_224 ( .gnd(gnd), .vdd(vdd), .A(_10308_), .B(_10149_), .Y(_10309_) );
NOR2X1 NOR2X1_815 ( .gnd(gnd), .vdd(vdd), .A(_10149_), .B(_10308_), .Y(_10310_) );
NOR2X1 NOR2X1_816 ( .gnd(gnd), .vdd(vdd), .A(_10310_), .B(_10309_), .Y(_10311_) );
OR2X2 OR2X2_241 ( .gnd(gnd), .vdd(vdd), .A(_10311_), .B(module_2_W_235_), .Y(_10312_) );
NAND2X1 NAND2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_235_), .B(_10311_), .Y(_10313_) );
NAND3X1 NAND3X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_10130_), .B(_10313_), .C(_10312_), .Y(_10314_) );
INVX2 INVX2_370 ( .gnd(gnd), .vdd(vdd), .A(_10314_), .Y(_10315_) );
AOI21X1 AOI21X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_10313_), .B(_10312_), .C(_10130_), .Y(_10316_) );
OAI21X1 OAI21X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_10315_), .B(_10316_), .C(_10148_), .Y(_10317_) );
INVX1 INVX1_1425 ( .gnd(gnd), .vdd(vdd), .A(_10317_), .Y(_10318_) );
OAI21X1 OAI21X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_10134_), .B(_9200_), .C(_10129_), .Y(_10319_) );
NOR2X1 NOR2X1_817 ( .gnd(gnd), .vdd(vdd), .A(_10316_), .B(_10315_), .Y(_10320_) );
AND2X2 AND2X2_225 ( .gnd(gnd), .vdd(vdd), .A(_10320_), .B(_10319_), .Y(_10321_) );
NOR2X1 NOR2X1_818 ( .gnd(gnd), .vdd(vdd), .A(_10318_), .B(_10321_), .Y(_10322_) );
INVX2 INVX2_371 ( .gnd(gnd), .vdd(vdd), .A(_10322_), .Y(_10323_) );
INVX1 INVX1_1426 ( .gnd(gnd), .vdd(vdd), .A(_10311_), .Y(_10324_) );
AOI21X1 AOI21X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_10013_), .B(_10011_), .C(_10031_), .Y(_10325_) );
OAI21X1 OAI21X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_9977_), .B(_9975_), .C(_9968_), .Y(_10326_) );
INVX1 INVX1_1427 ( .gnd(gnd), .vdd(vdd), .A(_10326_), .Y(_10327_) );
OR2X2 OR2X2_242 ( .gnd(gnd), .vdd(vdd), .A(_10277_), .B(_10279_), .Y(_10328_) );
OAI21X1 OAI21X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_9931_), .B(_9928_), .C(module_2_W_167_), .Y(_10329_) );
INVX1 INVX1_1428 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_167_), .Y(_10330_) );
NAND3X1 NAND3X1_2319 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_166_), .B(_10330_), .C(_9926_), .Y(_10331_) );
OR2X2 OR2X2_243 ( .gnd(gnd), .vdd(vdd), .A(_10266_), .B(_10269_), .Y(_10332_) );
INVX1 INVX1_1429 ( .gnd(gnd), .vdd(vdd), .A(_9855_), .Y(_10333_) );
AOI21X1 AOI21X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_9576_), .B(_9823_), .C(_9826_), .Y(_10334_) );
INVX1 INVX1_1430 ( .gnd(gnd), .vdd(vdd), .A(_10334_), .Y(_10335_) );
NOR2X1 NOR2X1_819 ( .gnd(gnd), .vdd(vdd), .A(_10235_), .B(_10237_), .Y(_10336_) );
OAI21X1 OAI21X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_9784_), .B(_9786_), .C(_9779_), .Y(_10337_) );
NOR2X1 NOR2X1_820 ( .gnd(gnd), .vdd(vdd), .A(_10224_), .B(_10226_), .Y(_10338_) );
OAI21X1 OAI21X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_9742_), .B(_9744_), .C(_9737_), .Y(_10339_) );
NOR2X1 NOR2X1_821 ( .gnd(gnd), .vdd(vdd), .A(_10213_), .B(_10216_), .Y(_10340_) );
INVX1 INVX1_1431 ( .gnd(gnd), .vdd(vdd), .A(_10340_), .Y(_10341_) );
AOI21X1 AOI21X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_9702_), .B(_9582_), .C(_9705_), .Y(_10342_) );
AOI21X1 AOI21X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_9667_), .B(_9584_), .C(_9670_), .Y(_10343_) );
AOI21X1 AOI21X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_9587_), .B(_9629_), .C(_9633_), .Y(_10344_) );
INVX1 INVX1_1432 ( .gnd(gnd), .vdd(vdd), .A(_9604_), .Y(_10345_) );
NOR2X1 NOR2X1_822 ( .gnd(gnd), .vdd(vdd), .A(_10345_), .B(_9609_), .Y(_10346_) );
XNOR2X1 XNOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_7_), .B(module_2_W_23_), .Y(_10347_) );
XOR2X1 XOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_12285_), .B(_10347_), .Y(_10348_) );
XNOR2X1 XNOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .B(module_2_W_11_), .Y(_10349_) );
XNOR2X1 XNOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_10349_), .B(_10348_), .Y(_10350_) );
XNOR2X1 XNOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_10350_), .B(_9599_), .Y(_10351_) );
NAND2X1 NAND2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_12293_), .B(_12295_), .Y(_10352_) );
XNOR2X1 XNOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_10352_), .B(bloque_datos[7]), .Y(_10353_) );
NOR2X1 NOR2X1_823 ( .gnd(gnd), .vdd(vdd), .A(_10351_), .B(_10353_), .Y(_10354_) );
AND2X2 AND2X2_226 ( .gnd(gnd), .vdd(vdd), .A(_10353_), .B(_10351_), .Y(_10355_) );
NOR2X1 NOR2X1_824 ( .gnd(gnd), .vdd(vdd), .A(_10354_), .B(_10355_), .Y(_10356_) );
NOR2X1 NOR2X1_825 ( .gnd(gnd), .vdd(vdd), .A(_10346_), .B(_10356_), .Y(_10357_) );
AND2X2 AND2X2_227 ( .gnd(gnd), .vdd(vdd), .A(_10356_), .B(_10346_), .Y(_10358_) );
OAI21X1 OAI21X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_10358_), .B(_10357_), .C(_10182_), .Y(_10359_) );
OR2X2 OR2X2_244 ( .gnd(gnd), .vdd(vdd), .A(_10356_), .B(_10346_), .Y(_10360_) );
NAND2X1 NAND2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_10346_), .B(_10356_), .Y(_10361_) );
NAND3X1 NAND3X1_2320 ( .gnd(gnd), .vdd(vdd), .A(_10184_), .B(_10361_), .C(_10360_), .Y(_10362_) );
AND2X2 AND2X2_228 ( .gnd(gnd), .vdd(vdd), .A(_10362_), .B(_10359_), .Y(_10363_) );
AOI21X1 AOI21X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_9624_), .B(_9623_), .C(_9622_), .Y(_10364_) );
OAI21X1 OAI21X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_12312_), .B(_12307_), .C(bloque_datos_23_bF_buf3_), .Y(_10365_) );
NAND2X1 NAND2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_12309_), .B(_12308_), .Y(_10366_) );
OR2X2 OR2X2_245 ( .gnd(gnd), .vdd(vdd), .A(_10366_), .B(bloque_datos_23_bF_buf2_), .Y(_10367_) );
NAND3X1 NAND3X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_10365_), .B(_10364_), .C(_10367_), .Y(_10368_) );
INVX1 INVX1_1433 ( .gnd(gnd), .vdd(vdd), .A(_10365_), .Y(_10369_) );
NOR2X1 NOR2X1_826 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf1_), .B(_10366_), .Y(_10370_) );
OAI21X1 OAI21X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_10370_), .B(_10369_), .C(_9621_), .Y(_10371_) );
AOI21X1 AOI21X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_10368_), .B(_10371_), .C(_10363_), .Y(_10372_) );
NAND2X1 NAND2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_10359_), .B(_10362_), .Y(_10373_) );
NAND2X1 NAND2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_10371_), .B(_10368_), .Y(_10374_) );
NOR2X1 NOR2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_10373_), .B(_10374_), .Y(_10375_) );
OAI21X1 OAI21X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_10375_), .B(_10372_), .C(_10344_), .Y(_10376_) );
INVX1 INVX1_1434 ( .gnd(gnd), .vdd(vdd), .A(_10344_), .Y(_10377_) );
NOR3X1 NOR3X1_291 ( .gnd(gnd), .vdd(vdd), .A(_10370_), .B(_10369_), .C(_9621_), .Y(_10378_) );
AOI21X1 AOI21X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_10365_), .B(_10367_), .C(_10364_), .Y(_10379_) );
OAI21X1 OAI21X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_10378_), .B(_10379_), .C(_10373_), .Y(_10380_) );
NAND3X1 NAND3X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_10368_), .B(_10371_), .C(_10363_), .Y(_10381_) );
NAND3X1 NAND3X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_10380_), .B(_10381_), .C(_10377_), .Y(_10382_) );
NAND3X1 NAND3X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_10190_), .B(_10382_), .C(_10376_), .Y(_10383_) );
OAI21X1 OAI21X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_10375_), .B(_10372_), .C(_10377_), .Y(_10384_) );
NAND3X1 NAND3X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_10344_), .B(_10380_), .C(_10381_), .Y(_10385_) );
NAND3X1 NAND3X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_10195_), .B(_10385_), .C(_10384_), .Y(_10386_) );
NAND2X1 NAND2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_10386_), .B(_10383_), .Y(_10387_) );
NAND2X1 NAND2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_12326_), .B(_12325_), .Y(_10388_) );
XNOR2X1 XNOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_10388_), .B(bloque_datos[39]), .Y(_10389_) );
NOR2X1 NOR2X1_828 ( .gnd(gnd), .vdd(vdd), .A(_9659_), .B(_10389_), .Y(_10390_) );
AND2X2 AND2X2_229 ( .gnd(gnd), .vdd(vdd), .A(_10389_), .B(_9659_), .Y(_10391_) );
OAI21X1 OAI21X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_10391_), .B(_10390_), .C(_10387_), .Y(_10392_) );
AND2X2 AND2X2_230 ( .gnd(gnd), .vdd(vdd), .A(_10383_), .B(_10386_), .Y(_10393_) );
OR2X2 OR2X2_246 ( .gnd(gnd), .vdd(vdd), .A(_10389_), .B(_9659_), .Y(_10394_) );
NAND2X1 NAND2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_9659_), .B(_10389_), .Y(_10395_) );
NAND3X1 NAND3X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_10394_), .B(_10395_), .C(_10393_), .Y(_10396_) );
NAND3X1 NAND3X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_10343_), .B(_10392_), .C(_10396_), .Y(_10397_) );
OAI21X1 OAI21X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_9669_), .B(_9671_), .C(_9664_), .Y(_10398_) );
AOI21X1 AOI21X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_10394_), .B(_10395_), .C(_10393_), .Y(_10399_) );
NOR3X1 NOR3X1_292 ( .gnd(gnd), .vdd(vdd), .A(_10390_), .B(_10391_), .C(_10387_), .Y(_10400_) );
OAI21X1 OAI21X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_10399_), .B(_10400_), .C(_10398_), .Y(_10401_) );
NAND3X1 NAND3X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_10205_), .B(_10397_), .C(_10401_), .Y(_10402_) );
NAND3X1 NAND3X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_10398_), .B(_10392_), .C(_10396_), .Y(_10403_) );
OAI21X1 OAI21X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_10399_), .B(_10400_), .C(_10343_), .Y(_10404_) );
NAND3X1 NAND3X1_2331 ( .gnd(gnd), .vdd(vdd), .A(_10207_), .B(_10403_), .C(_10404_), .Y(_10405_) );
AND2X2 AND2X2_231 ( .gnd(gnd), .vdd(vdd), .A(_10402_), .B(_10405_), .Y(_10406_) );
XNOR2X1 XNOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_12335_), .B(bloque_datos[55]), .Y(_10407_) );
OR2X2 OR2X2_247 ( .gnd(gnd), .vdd(vdd), .A(_10407_), .B(_9694_), .Y(_10408_) );
NAND2X1 NAND2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_9694_), .B(_10407_), .Y(_10409_) );
AOI21X1 AOI21X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_10409_), .B(_10408_), .C(_10406_), .Y(_10410_) );
NAND2X1 NAND2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_10402_), .B(_10405_), .Y(_10411_) );
NOR2X1 NOR2X1_829 ( .gnd(gnd), .vdd(vdd), .A(_9694_), .B(_10407_), .Y(_10412_) );
AND2X2 AND2X2_232 ( .gnd(gnd), .vdd(vdd), .A(_10407_), .B(_9694_), .Y(_10413_) );
NOR3X1 NOR3X1_293 ( .gnd(gnd), .vdd(vdd), .A(_10413_), .B(_10412_), .C(_10411_), .Y(_10414_) );
OAI21X1 OAI21X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_10410_), .B(_10414_), .C(_10342_), .Y(_10415_) );
OAI21X1 OAI21X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_9704_), .B(_9706_), .C(_9699_), .Y(_10416_) );
OAI21X1 OAI21X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_10413_), .B(_10412_), .C(_10411_), .Y(_10417_) );
NAND3X1 NAND3X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_10409_), .B(_10408_), .C(_10406_), .Y(_10418_) );
NAND3X1 NAND3X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_10417_), .B(_10416_), .C(_10418_), .Y(_10419_) );
NAND3X1 NAND3X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_10341_), .B(_10419_), .C(_10415_), .Y(_10420_) );
OAI21X1 OAI21X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_10410_), .B(_10414_), .C(_10416_), .Y(_10421_) );
NAND3X1 NAND3X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_10342_), .B(_10417_), .C(_10418_), .Y(_10422_) );
NAND3X1 NAND3X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_10340_), .B(_10422_), .C(_10421_), .Y(_10423_) );
AND2X2 AND2X2_233 ( .gnd(gnd), .vdd(vdd), .A(_10420_), .B(_10423_), .Y(_10424_) );
OAI21X1 OAI21X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_12341_), .B(_12347_), .C(bloque_datos_71_bF_buf3_), .Y(_10425_) );
INVX1 INVX1_1435 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf2_), .Y(_10426_) );
OAI21X1 OAI21X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_12343_), .B(_12346_), .C(_12342_), .Y(_10427_) );
NAND3X1 NAND3X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_12272_), .B(_12340_), .C(_12337_), .Y(_10428_) );
NAND3X1 NAND3X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_10426_), .B(_10427_), .C(_10428_), .Y(_10429_) );
NAND2X1 NAND2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_10429_), .B(_10425_), .Y(_10430_) );
OR2X2 OR2X2_248 ( .gnd(gnd), .vdd(vdd), .A(_10430_), .B(_9732_), .Y(_10431_) );
NAND2X1 NAND2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_9732_), .B(_10430_), .Y(_10432_) );
AOI21X1 AOI21X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_10431_), .B(_10432_), .C(_10424_), .Y(_10433_) );
NAND2X1 NAND2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_10420_), .B(_10423_), .Y(_10434_) );
NOR2X1 NOR2X1_830 ( .gnd(gnd), .vdd(vdd), .A(_9732_), .B(_10430_), .Y(_10435_) );
AND2X2 AND2X2_234 ( .gnd(gnd), .vdd(vdd), .A(_10430_), .B(_9732_), .Y(_10436_) );
NOR3X1 NOR3X1_294 ( .gnd(gnd), .vdd(vdd), .A(_10436_), .B(_10435_), .C(_10434_), .Y(_10437_) );
OAI21X1 OAI21X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_10433_), .B(_10437_), .C(_10339_), .Y(_10438_) );
AOI21X1 AOI21X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_9740_), .B(_9580_), .C(_9743_), .Y(_10439_) );
OAI21X1 OAI21X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_10436_), .B(_10435_), .C(_10434_), .Y(_10440_) );
NAND3X1 NAND3X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_10431_), .B(_10432_), .C(_10424_), .Y(_10441_) );
NAND3X1 NAND3X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_10439_), .B(_10440_), .C(_10441_), .Y(_10442_) );
AOI21X1 AOI21X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_10442_), .B(_10438_), .C(_10338_), .Y(_10443_) );
INVX1 INVX1_1436 ( .gnd(gnd), .vdd(vdd), .A(_10338_), .Y(_10444_) );
OAI21X1 OAI21X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_10433_), .B(_10437_), .C(_10439_), .Y(_10445_) );
NAND3X1 NAND3X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_10440_), .B(_10339_), .C(_10441_), .Y(_10446_) );
AOI21X1 AOI21X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_10446_), .B(_10445_), .C(_10444_), .Y(_10447_) );
OR2X2 OR2X2_249 ( .gnd(gnd), .vdd(vdd), .A(_10443_), .B(_10447_), .Y(_10448_) );
NAND3X1 NAND3X1_2342 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf1_), .B(_12357_), .C(_12361_), .Y(_10449_) );
INVX1 INVX1_1437 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf0_), .Y(_10450_) );
OAI21X1 OAI21X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_12358_), .B(_12356_), .C(_10450_), .Y(_10451_) );
NAND2X1 NAND2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_10449_), .B(_10451_), .Y(_10452_) );
OR2X2 OR2X2_250 ( .gnd(gnd), .vdd(vdd), .A(_10452_), .B(_9774_), .Y(_10453_) );
NAND2X1 NAND2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_9774_), .B(_10452_), .Y(_10454_) );
NAND3X1 NAND3X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_10453_), .B(_10454_), .C(_10448_), .Y(_10455_) );
NOR2X1 NOR2X1_831 ( .gnd(gnd), .vdd(vdd), .A(_10443_), .B(_10447_), .Y(_10456_) );
NOR2X1 NOR2X1_832 ( .gnd(gnd), .vdd(vdd), .A(_9774_), .B(_10452_), .Y(_10457_) );
AND2X2 AND2X2_235 ( .gnd(gnd), .vdd(vdd), .A(_10452_), .B(_9774_), .Y(_10458_) );
OAI21X1 OAI21X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_10458_), .B(_10457_), .C(_10456_), .Y(_10459_) );
NAND3X1 NAND3X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_10459_), .B(_10337_), .C(_10455_), .Y(_10460_) );
AOI21X1 AOI21X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_9782_), .B(_9578_), .C(_9785_), .Y(_10461_) );
NOR3X1 NOR3X1_295 ( .gnd(gnd), .vdd(vdd), .A(_10458_), .B(_10457_), .C(_10456_), .Y(_10462_) );
AOI21X1 AOI21X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_10454_), .B(_10453_), .C(_10448_), .Y(_10463_) );
OAI21X1 OAI21X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_10462_), .B(_10463_), .C(_10461_), .Y(_10464_) );
AOI21X1 AOI21X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_10460_), .B(_10464_), .C(_10336_), .Y(_10465_) );
INVX1 INVX1_1438 ( .gnd(gnd), .vdd(vdd), .A(_10336_), .Y(_10466_) );
NAND3X1 NAND3X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_10461_), .B(_10459_), .C(_10455_), .Y(_10467_) );
OAI21X1 OAI21X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_10462_), .B(_10463_), .C(_10337_), .Y(_10468_) );
AOI21X1 AOI21X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_10467_), .B(_10468_), .C(_10466_), .Y(_10469_) );
NOR2X1 NOR2X1_833 ( .gnd(gnd), .vdd(vdd), .A(_10465_), .B(_10469_), .Y(_10470_) );
NAND3X1 NAND3X1_2346 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_135_), .B(_12369_), .C(_12372_), .Y(_10471_) );
INVX1 INVX1_1439 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_135_), .Y(_10472_) );
OAI21X1 OAI21X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_12370_), .B(_12368_), .C(_10472_), .Y(_10473_) );
NAND2X1 NAND2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_10471_), .B(_10473_), .Y(_10474_) );
NOR2X1 NOR2X1_834 ( .gnd(gnd), .vdd(vdd), .A(_10474_), .B(_9815_), .Y(_10475_) );
NAND2X1 NAND2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_10474_), .B(_9815_), .Y(_10476_) );
INVX1 INVX1_1440 ( .gnd(gnd), .vdd(vdd), .A(_10476_), .Y(_10477_) );
NOR3X1 NOR3X1_296 ( .gnd(gnd), .vdd(vdd), .A(_10477_), .B(_10475_), .C(_10470_), .Y(_10478_) );
OR2X2 OR2X2_251 ( .gnd(gnd), .vdd(vdd), .A(_10465_), .B(_10469_), .Y(_10479_) );
INVX1 INVX1_1441 ( .gnd(gnd), .vdd(vdd), .A(_10475_), .Y(_10480_) );
AOI21X1 AOI21X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_10476_), .B(_10480_), .C(_10479_), .Y(_10481_) );
OAI21X1 OAI21X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_10478_), .B(_10481_), .C(_10335_), .Y(_10482_) );
NAND3X1 NAND3X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_10476_), .B(_10480_), .C(_10479_), .Y(_10483_) );
OAI21X1 OAI21X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_10477_), .B(_10475_), .C(_10470_), .Y(_10484_) );
NAND3X1 NAND3X1_2348 ( .gnd(gnd), .vdd(vdd), .A(_10334_), .B(_10484_), .C(_10483_), .Y(_10485_) );
AOI21X1 AOI21X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_10485_), .B(_10482_), .C(_10249_), .Y(_10486_) );
INVX1 INVX1_1442 ( .gnd(gnd), .vdd(vdd), .A(_10249_), .Y(_10487_) );
OAI21X1 OAI21X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_10478_), .B(_10481_), .C(_10334_), .Y(_10488_) );
NAND3X1 NAND3X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_10484_), .B(_10483_), .C(_10335_), .Y(_10489_) );
AOI21X1 AOI21X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_10489_), .B(_10488_), .C(_10487_), .Y(_10490_) );
OAI21X1 OAI21X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_10486_), .B(_10490_), .C(_10333_), .Y(_10491_) );
NAND3X1 NAND3X1_2350 ( .gnd(gnd), .vdd(vdd), .A(_10487_), .B(_10489_), .C(_10488_), .Y(_10492_) );
NAND3X1 NAND3X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_10249_), .B(_10485_), .C(_10482_), .Y(_10493_) );
NAND3X1 NAND3X1_2352 ( .gnd(gnd), .vdd(vdd), .A(_9855_), .B(_10492_), .C(_10493_), .Y(_10494_) );
NAND2X1 NAND2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_10494_), .B(_10491_), .Y(_10495_) );
OAI21X1 OAI21X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_9866_), .B(_9888_), .C(_10495_), .Y(_10496_) );
INVX1 INVX1_1443 ( .gnd(gnd), .vdd(vdd), .A(_12381_), .Y(_10497_) );
OAI21X1 OAI21X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_9865_), .B(_9867_), .C(_9860_), .Y(_10498_) );
INVX1 INVX1_1444 ( .gnd(gnd), .vdd(vdd), .A(_10498_), .Y(_10499_) );
AND2X2 AND2X2_236 ( .gnd(gnd), .vdd(vdd), .A(_10491_), .B(_10494_), .Y(_10500_) );
AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_12378_), .B(_10497_), .C(_10500_), .D(_10499_), .Y(_10501_) );
NAND3X1 NAND3X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_10258_), .B(_10496_), .C(_10501_), .Y(_10502_) );
INVX1 INVX1_1445 ( .gnd(gnd), .vdd(vdd), .A(_10258_), .Y(_10503_) );
NOR2X1 NOR2X1_835 ( .gnd(gnd), .vdd(vdd), .A(_10499_), .B(_10500_), .Y(_10504_) );
NAND2X1 NAND2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_12378_), .B(_10497_), .Y(_10505_) );
OAI21X1 OAI21X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_10495_), .B(_10498_), .C(_10505_), .Y(_10506_) );
OAI21X1 OAI21X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_10504_), .B(_10506_), .C(_10503_), .Y(_10507_) );
AND2X2 AND2X2_237 ( .gnd(gnd), .vdd(vdd), .A(_10502_), .B(_10507_), .Y(_10508_) );
INVX1 INVX1_1446 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_151_), .Y(_10509_) );
AOI21X1 AOI21X1_1463 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_150_), .B(_9891_), .C(_10509_), .Y(_10510_) );
NOR3X1 NOR3X1_297 ( .gnd(gnd), .vdd(vdd), .A(_9893_), .B(module_2_W_151_), .C(_9896_), .Y(_10511_) );
OAI21X1 OAI21X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_10510_), .B(_10511_), .C(_10508_), .Y(_10512_) );
NAND2X1 NAND2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_10507_), .B(_10502_), .Y(_10513_) );
OAI21X1 OAI21X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_9896_), .B(_9893_), .C(module_2_W_151_), .Y(_10514_) );
NAND3X1 NAND3X1_2354 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_150_), .B(_10509_), .C(_9891_), .Y(_10515_) );
NAND3X1 NAND3X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_10514_), .B(_10515_), .C(_10513_), .Y(_10516_) );
AND2X2 AND2X2_238 ( .gnd(gnd), .vdd(vdd), .A(_10512_), .B(_10516_), .Y(_10517_) );
OAI21X1 OAI21X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_9922_), .B(_9902_), .C(_10517_), .Y(_10518_) );
OAI21X1 OAI21X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_9570_), .B(_9923_), .C(_9905_), .Y(_10519_) );
INVX1 INVX1_1447 ( .gnd(gnd), .vdd(vdd), .A(_10519_), .Y(_10520_) );
NAND2X1 NAND2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_10516_), .B(_10512_), .Y(_10521_) );
AOI21X1 AOI21X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_10521_), .B(_10520_), .C(_12393_), .Y(_10522_) );
NAND3X1 NAND3X1_2356 ( .gnd(gnd), .vdd(vdd), .A(_10332_), .B(_10518_), .C(_10522_), .Y(_10523_) );
NOR2X1 NOR2X1_836 ( .gnd(gnd), .vdd(vdd), .A(_10521_), .B(_10520_), .Y(_10524_) );
INVX1 INVX1_1448 ( .gnd(gnd), .vdd(vdd), .A(_12393_), .Y(_10525_) );
OAI21X1 OAI21X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_10517_), .B(_10519_), .C(_10525_), .Y(_10526_) );
OAI21X1 OAI21X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_10526_), .B(_10524_), .C(_10271_), .Y(_10527_) );
NAND2X1 NAND2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_10523_), .B(_10527_), .Y(_10528_) );
AOI21X1 AOI21X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_10329_), .B(_10331_), .C(_10528_), .Y(_10529_) );
NAND3X1 NAND3X1_2357 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_166_), .B(module_2_W_167_), .C(_9926_), .Y(_10530_) );
OAI21X1 OAI21X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_9931_), .B(_9928_), .C(_10330_), .Y(_10531_) );
AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_10523_), .B(_10527_), .C(_10531_), .D(_10530_), .Y(_10532_) );
NOR2X1 NOR2X1_837 ( .gnd(gnd), .vdd(vdd), .A(_10532_), .B(_10529_), .Y(_10533_) );
OAI21X1 OAI21X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_9957_), .B(_9937_), .C(_10533_), .Y(_10534_) );
OAI21X1 OAI21X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_9958_), .B(_9568_), .C(_9940_), .Y(_10535_) );
INVX1 INVX1_1449 ( .gnd(gnd), .vdd(vdd), .A(_10535_), .Y(_10536_) );
NAND2X1 NAND2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_10530_), .B(_10531_), .Y(_10537_) );
XNOR2X1 XNOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_10537_), .B(_10528_), .Y(_10538_) );
AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_12401_), .B(_12403_), .C(_10538_), .D(_10536_), .Y(_10539_) );
NAND3X1 NAND3X1_2358 ( .gnd(gnd), .vdd(vdd), .A(_10328_), .B(_10534_), .C(_10539_), .Y(_10540_) );
NOR2X1 NOR2X1_838 ( .gnd(gnd), .vdd(vdd), .A(_10538_), .B(_10536_), .Y(_10541_) );
OAI21X1 OAI21X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_10533_), .B(_10535_), .C(_12404_), .Y(_10542_) );
OAI21X1 OAI21X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_10541_), .B(_10542_), .C(_10281_), .Y(_10543_) );
AND2X2 AND2X2_239 ( .gnd(gnd), .vdd(vdd), .A(_10540_), .B(_10543_), .Y(_10544_) );
INVX1 INVX1_1450 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_183_), .Y(_10545_) );
AOI21X1 AOI21X1_1466 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_182_), .B(_9961_), .C(_10545_), .Y(_10546_) );
NOR3X1 NOR3X1_298 ( .gnd(gnd), .vdd(vdd), .A(_9963_), .B(module_2_W_183_), .C(_9966_), .Y(_10547_) );
OAI21X1 OAI21X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_10546_), .B(_10547_), .C(_10544_), .Y(_10548_) );
NAND2X1 NAND2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_10543_), .B(_10540_), .Y(_10549_) );
OAI21X1 OAI21X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_9966_), .B(_9963_), .C(module_2_W_183_), .Y(_10550_) );
NAND3X1 NAND3X1_2359 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_182_), .B(_10545_), .C(_9961_), .Y(_10551_) );
NAND3X1 NAND3X1_2360 ( .gnd(gnd), .vdd(vdd), .A(_10550_), .B(_10551_), .C(_10549_), .Y(_10552_) );
NAND2X1 NAND2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_10552_), .B(_10548_), .Y(_10553_) );
NOR2X1 NOR2X1_839 ( .gnd(gnd), .vdd(vdd), .A(_10553_), .B(_10327_), .Y(_10554_) );
AND2X2 AND2X2_240 ( .gnd(gnd), .vdd(vdd), .A(_10548_), .B(_10552_), .Y(_10555_) );
OAI21X1 OAI21X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_10555_), .B(_10326_), .C(_8986_), .Y(_10556_) );
OAI21X1 OAI21X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_10556_), .B(_10554_), .C(module_2_W_199_), .Y(_10557_) );
INVX1 INVX1_1451 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_199_), .Y(_10558_) );
OAI21X1 OAI21X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_9976_), .B(_9995_), .C(_10555_), .Y(_10560_) );
AOI21X1 AOI21X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_10553_), .B(_10327_), .C(_12418_), .Y(_10561_) );
NAND3X1 NAND3X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_10558_), .B(_10560_), .C(_10561_), .Y(_10562_) );
NAND2X1 NAND2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_10562_), .B(_10557_), .Y(_10563_) );
NOR3X1 NOR3X1_299 ( .gnd(gnd), .vdd(vdd), .A(_9995_), .B(_9997_), .C(_9996_), .Y(_10564_) );
NOR3X1 NOR3X1_300 ( .gnd(gnd), .vdd(vdd), .A(_9562_), .B(_10002_), .C(_10564_), .Y(_10565_) );
OAI21X1 OAI21X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_10565_), .B(_10001_), .C(_10290_), .Y(_10566_) );
INVX2 INVX2_372 ( .gnd(gnd), .vdd(vdd), .A(_10290_), .Y(_10567_) );
NAND3X1 NAND3X1_2362 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_198_), .B(_10567_), .C(_9999_), .Y(_10568_) );
NAND3X1 NAND3X1_2363 ( .gnd(gnd), .vdd(vdd), .A(_10566_), .B(_10568_), .C(_10563_), .Y(_10569_) );
AND2X2 AND2X2_241 ( .gnd(gnd), .vdd(vdd), .A(_10557_), .B(_10562_), .Y(_10571_) );
AOI21X1 AOI21X1_1468 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_198_), .B(_9999_), .C(_10567_), .Y(_10572_) );
INVX1 INVX1_1452 ( .gnd(gnd), .vdd(vdd), .A(_10568_), .Y(_10573_) );
OAI21X1 OAI21X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_10573_), .B(_10572_), .C(_10571_), .Y(_10574_) );
AOI21X1 AOI21X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_10569_), .B(_10574_), .C(_10325_), .Y(_10575_) );
OAI21X1 OAI21X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_10032_), .B(_9561_), .C(_10012_), .Y(_10576_) );
NAND2X1 NAND2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_10569_), .B(_10574_), .Y(_10577_) );
OAI21X1 OAI21X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_10577_), .B(_10576_), .C(_12433_), .Y(_10578_) );
NOR3X1 NOR3X1_301 ( .gnd(gnd), .vdd(vdd), .A(_10575_), .B(_10301_), .C(_10578_), .Y(_10579_) );
INVX2 INVX2_373 ( .gnd(gnd), .vdd(vdd), .A(_10301_), .Y(_10580_) );
INVX1 INVX1_1453 ( .gnd(gnd), .vdd(vdd), .A(_10575_), .Y(_10582_) );
AND2X2 AND2X2_242 ( .gnd(gnd), .vdd(vdd), .A(_10574_), .B(_10569_), .Y(_10583_) );
AOI21X1 AOI21X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_10325_), .B(_10583_), .C(_12436_), .Y(_10584_) );
AOI21X1 AOI21X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_10582_), .B(_10584_), .C(_10580_), .Y(_10585_) );
NOR2X1 NOR2X1_840 ( .gnd(gnd), .vdd(vdd), .A(_10579_), .B(_10585_), .Y(_10586_) );
INVX1 INVX1_1454 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_215_), .Y(_10587_) );
AOI21X1 AOI21X1_1472 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_214_), .B(_10035_), .C(_10587_), .Y(_10588_) );
NOR3X1 NOR3X1_302 ( .gnd(gnd), .vdd(vdd), .A(_10037_), .B(module_2_W_215_), .C(_10040_), .Y(_10589_) );
OAI21X1 OAI21X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_10588_), .B(_10589_), .C(_10586_), .Y(_10590_) );
NAND3X1 NAND3X1_2364 ( .gnd(gnd), .vdd(vdd), .A(_10580_), .B(_10582_), .C(_10584_), .Y(_10591_) );
OAI21X1 OAI21X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_10578_), .B(_10575_), .C(_10301_), .Y(_10593_) );
NAND2X1 NAND2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_10593_), .B(_10591_), .Y(_10594_) );
OAI21X1 OAI21X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_10040_), .B(_10037_), .C(module_2_W_215_), .Y(_10595_) );
NAND3X1 NAND3X1_2365 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_214_), .B(_10587_), .C(_10035_), .Y(_10596_) );
NAND3X1 NAND3X1_2366 ( .gnd(gnd), .vdd(vdd), .A(_10595_), .B(_10596_), .C(_10594_), .Y(_10597_) );
AND2X2 AND2X2_243 ( .gnd(gnd), .vdd(vdd), .A(_10590_), .B(_10597_), .Y(_10598_) );
OAI21X1 OAI21X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_10068_), .B(_10046_), .C(_10598_), .Y(_10599_) );
AOI21X1 AOI21X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_10050_), .B(_10048_), .C(_10068_), .Y(_10600_) );
NAND2X1 NAND2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_10597_), .B(_10590_), .Y(_10601_) );
AOI21X1 AOI21X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_10600_), .B(_10601_), .C(_12445_), .Y(_10602_) );
NAND3X1 NAND3X1_2367 ( .gnd(gnd), .vdd(vdd), .A(_10324_), .B(_10602_), .C(_10599_), .Y(_10604_) );
NOR2X1 NOR2X1_841 ( .gnd(gnd), .vdd(vdd), .A(_10600_), .B(_10601_), .Y(_10605_) );
INVX1 INVX1_1455 ( .gnd(gnd), .vdd(vdd), .A(_12445_), .Y(_10606_) );
OAI21X1 OAI21X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_10069_), .B(_9558_), .C(_10049_), .Y(_10607_) );
OAI21X1 OAI21X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_10598_), .B(_10607_), .C(_10606_), .Y(_10608_) );
OAI21X1 OAI21X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_10608_), .B(_10605_), .C(_10311_), .Y(_10609_) );
AND2X2 AND2X2_244 ( .gnd(gnd), .vdd(vdd), .A(_10609_), .B(_10604_), .Y(_10610_) );
INVX1 INVX1_1456 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_231_), .Y(_10611_) );
AOI21X1 AOI21X1_1475 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_230_), .B(_10072_), .C(_10611_), .Y(_10612_) );
NOR3X1 NOR3X1_303 ( .gnd(gnd), .vdd(vdd), .A(_10074_), .B(module_2_W_231_), .C(_10077_), .Y(_10613_) );
OAI21X1 OAI21X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_10612_), .B(_10613_), .C(_10610_), .Y(_10615_) );
NAND2X1 NAND2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_10604_), .B(_10609_), .Y(_10616_) );
OAI21X1 OAI21X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_10077_), .B(_10074_), .C(module_2_W_231_), .Y(_10617_) );
NAND3X1 NAND3X1_2368 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_230_), .B(_10611_), .C(_10072_), .Y(_10618_) );
NAND3X1 NAND3X1_2369 ( .gnd(gnd), .vdd(vdd), .A(_10617_), .B(_10618_), .C(_10616_), .Y(_10619_) );
AND2X2 AND2X2_245 ( .gnd(gnd), .vdd(vdd), .A(_10615_), .B(_10619_), .Y(_10620_) );
OAI21X1 OAI21X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_10105_), .B(_10083_), .C(_10620_), .Y(_10621_) );
OAI21X1 OAI21X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_10106_), .B(_9552_), .C(_10086_), .Y(_10622_) );
INVX1 INVX1_1457 ( .gnd(gnd), .vdd(vdd), .A(_10622_), .Y(_10623_) );
NAND2X1 NAND2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_10619_), .B(_10615_), .Y(_10624_) );
AOI21X1 AOI21X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_10624_), .B(_10623_), .C(_12458_), .Y(_10626_) );
NAND3X1 NAND3X1_2370 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_247_), .B(_10621_), .C(_10626_), .Y(_10627_) );
INVX2 INVX2_374 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_247_), .Y(_10628_) );
NOR2X1 NOR2X1_842 ( .gnd(gnd), .vdd(vdd), .A(_10624_), .B(_10623_), .Y(_10629_) );
INVX1 INVX1_1458 ( .gnd(gnd), .vdd(vdd), .A(_12458_), .Y(_10630_) );
OAI21X1 OAI21X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_10620_), .B(_10622_), .C(_10630_), .Y(_10631_) );
OAI21X1 OAI21X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_10631_), .B(_10629_), .C(_10628_), .Y(_10632_) );
NAND3X1 NAND3X1_2371 ( .gnd(gnd), .vdd(vdd), .A(_10627_), .B(_10632_), .C(_10110_), .Y(_10633_) );
NOR2X1 NOR2X1_843 ( .gnd(gnd), .vdd(vdd), .A(_10111_), .B(_10114_), .Y(_10634_) );
NOR3X1 NOR3X1_304 ( .gnd(gnd), .vdd(vdd), .A(_10629_), .B(_10628_), .C(_10631_), .Y(_10635_) );
AOI21X1 AOI21X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_10621_), .B(_10626_), .C(module_2_W_247_), .Y(_10637_) );
OAI21X1 OAI21X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_10635_), .B(_10637_), .C(_10634_), .Y(_10638_) );
NAND3X1 NAND3X1_2372 ( .gnd(gnd), .vdd(vdd), .A(_10323_), .B(_10633_), .C(_10638_), .Y(_10639_) );
NAND3X1 NAND3X1_2373 ( .gnd(gnd), .vdd(vdd), .A(_10628_), .B(_10621_), .C(_10626_), .Y(_10640_) );
OAI21X1 OAI21X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_10631_), .B(_10629_), .C(module_2_W_247_), .Y(_10641_) );
AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_246_), .B(_10109_), .C(_10641_), .D(_10640_), .Y(_10642_) );
AOI21X1 AOI21X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_10627_), .B(_10632_), .C(_10110_), .Y(_10643_) );
OAI21X1 OAI21X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_10643_), .B(_10642_), .C(_10322_), .Y(_10644_) );
NAND3X1 NAND3X1_2374 ( .gnd(gnd), .vdd(vdd), .A(_10639_), .B(_10644_), .C(_10147_), .Y(_10645_) );
AOI21X1 AOI21X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_10110_), .B(_10115_), .C(_9527_), .Y(_10646_) );
OAI21X1 OAI21X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_10646_), .B(_9550_), .C(_10122_), .Y(_10648_) );
NOR3X1 NOR3X1_305 ( .gnd(gnd), .vdd(vdd), .A(_10642_), .B(_10322_), .C(_10643_), .Y(_10649_) );
AOI21X1 AOI21X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_10638_), .C(_10323_), .Y(_10650_) );
OAI21X1 OAI21X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_10649_), .B(_10650_), .C(_10648_), .Y(_10651_) );
NAND2X1 NAND2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_10651_), .B(_10645_), .Y(_10652_) );
NAND2X1 NAND2X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_10652_), .B(_10145_), .Y(_10653_) );
OAI21X1 OAI21X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_10649_), .B(_10650_), .C(_10147_), .Y(_10654_) );
NAND3X1 NAND3X1_2375 ( .gnd(gnd), .vdd(vdd), .A(_10639_), .B(_10644_), .C(_10648_), .Y(_10655_) );
NAND2X1 NAND2X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_10655_), .B(_10654_), .Y(_10656_) );
NAND3X1 NAND3X1_2376 ( .gnd(gnd), .vdd(vdd), .A(_9549_), .B(_10656_), .C(_10142_), .Y(_10657_) );
NAND2X1 NAND2X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_10657_), .B(_10653_), .Y(module_2_H_7_) );
NOR2X1 NOR2X1_844 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_248_), .B(_9074_), .Y(_10659_) );
INVX1 INVX1_1459 ( .gnd(gnd), .vdd(vdd), .A(_10659_), .Y(_10660_) );
OAI21X1 OAI21X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_9069_), .B(_9068_), .C(module_2_W_248_), .Y(_10661_) );
NAND2X1 NAND2X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_10661_), .B(_10660_), .Y(module_2_H_16_) );
XNOR2X1 XNOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_9201_), .B(module_2_W_249_), .Y(_10662_) );
INVX1 INVX1_1460 ( .gnd(gnd), .vdd(vdd), .A(_10662_), .Y(_10663_) );
OAI21X1 OAI21X1_1687 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_248_), .B(_9074_), .C(_10663_), .Y(_10664_) );
INVX2 INVX2_375 ( .gnd(gnd), .vdd(vdd), .A(_10664_), .Y(_10665_) );
NOR2X1 NOR2X1_845 ( .gnd(gnd), .vdd(vdd), .A(_10660_), .B(_10663_), .Y(_10666_) );
NOR2X1 NOR2X1_846 ( .gnd(gnd), .vdd(vdd), .A(_10666_), .B(_10665_), .Y(module_2_H_17_) );
NOR2X1 NOR2X1_847 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_249_), .B(_9544_), .Y(_10668_) );
INVX1 INVX1_1461 ( .gnd(gnd), .vdd(vdd), .A(_10668_), .Y(_10669_) );
NAND2X1 NAND2X1_1407 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_250_), .B(_10136_), .Y(_10670_) );
OR2X2 OR2X2_252 ( .gnd(gnd), .vdd(vdd), .A(_10136_), .B(module_2_W_250_), .Y(_10671_) );
AOI21X1 AOI21X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_10670_), .B(_10671_), .C(_10669_), .Y(_10672_) );
INVX1 INVX1_1462 ( .gnd(gnd), .vdd(vdd), .A(_10672_), .Y(_10673_) );
NAND3X1 NAND3X1_2377 ( .gnd(gnd), .vdd(vdd), .A(_10669_), .B(_10670_), .C(_10671_), .Y(_10674_) );
NAND2X1 NAND2X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_10674_), .B(_10673_), .Y(_10675_) );
XNOR2X1 XNOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_10675_), .B(_10665_), .Y(module_2_H_18_) );
OAI21X1 OAI21X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_10672_), .B(_10664_), .C(_10674_), .Y(_10677_) );
NOR2X1 NOR2X1_848 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_250_), .B(_10137_), .Y(_10678_) );
INVX1 INVX1_1463 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_251_), .Y(_10679_) );
OAI21X1 OAI21X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_10321_), .B(_10318_), .C(_10679_), .Y(_10680_) );
NAND2X1 NAND2X1_1409 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_251_), .B(_10322_), .Y(_10681_) );
NAND3X1 NAND3X1_2378 ( .gnd(gnd), .vdd(vdd), .A(_10678_), .B(_10680_), .C(_10681_), .Y(_10682_) );
AOI21X1 AOI21X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_10680_), .B(_10681_), .C(_10678_), .Y(_10683_) );
INVX1 INVX1_1464 ( .gnd(gnd), .vdd(vdd), .A(_10683_), .Y(_10684_) );
NAND2X1 NAND2X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_10682_), .B(_10684_), .Y(_10685_) );
XNOR2X1 XNOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_10685_), .B(_10677_), .Y(module_2_H_19_) );
AOI21X1 AOI21X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_10677_), .B(_10682_), .C(_10683_), .Y(_10687_) );
OAI21X1 OAI21X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .B(_10316_), .C(_10314_), .Y(_10688_) );
INVX2 INVX2_376 ( .gnd(gnd), .vdd(vdd), .A(_10313_), .Y(_10689_) );
OAI21X1 OAI21X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_10303_), .B(_10302_), .C(_10093_), .Y(_10690_) );
AOI21X1 AOI21X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_10690_), .B(_10149_), .C(_10304_), .Y(_10691_) );
NOR3X1 NOR3X1_306 ( .gnd(gnd), .vdd(vdd), .A(_10056_), .B(_10292_), .C(_10295_), .Y(_10692_) );
AOI21X1 AOI21X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_10296_), .B(_10299_), .C(_10692_), .Y(_10693_) );
OAI21X1 OAI21X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_10288_), .B(_10285_), .C(_10283_), .Y(_10694_) );
INVX1 INVX1_1465 ( .gnd(gnd), .vdd(vdd), .A(_10282_), .Y(_10695_) );
OR2X2 OR2X2_253 ( .gnd(gnd), .vdd(vdd), .A(_10273_), .B(_10156_), .Y(_10696_) );
OAI21X1 OAI21X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_10275_), .B(_10154_), .C(_10696_), .Y(_10698_) );
NOR2X1 NOR2X1_849 ( .gnd(gnd), .vdd(vdd), .A(_10157_), .B(_10332_), .Y(_10699_) );
OAI21X1 OAI21X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_10260_), .B(_10261_), .C(_9946_), .Y(_10700_) );
AOI21X1 AOI21X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_10700_), .B(_10158_), .C(_10262_), .Y(_10701_) );
OAI21X1 OAI21X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_10256_), .B(_10160_), .C(_10252_), .Y(_10702_) );
INVX2 INVX2_377 ( .gnd(gnd), .vdd(vdd), .A(_10702_), .Y(_10703_) );
NAND2X1 NAND2X1_1411 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_139_), .B(_10249_), .Y(_10704_) );
AND2X2 AND2X2_246 ( .gnd(gnd), .vdd(vdd), .A(_10246_), .B(_10242_), .Y(_10705_) );
INVX1 INVX1_1466 ( .gnd(gnd), .vdd(vdd), .A(_10243_), .Y(_10706_) );
INVX1 INVX1_1467 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf3_), .Y(_10707_) );
XNOR2X1 XNOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_8878_), .B(_11202_), .Y(_10709_) );
NAND2X1 NAND2X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_10231_), .B(_10236_), .Y(_10710_) );
XOR2X1 XOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_8853_), .B(_10730_), .Y(_10711_) );
INVX1 INVX1_1468 ( .gnd(gnd), .vdd(vdd), .A(_10165_), .Y(_10712_) );
AOI21X1 AOI21X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_10219_), .B(_10217_), .C(_9793_), .Y(_10713_) );
OAI21X1 OAI21X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_10712_), .B(_10713_), .C(_10220_), .Y(_10714_) );
XNOR2X1 XNOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_8827_), .B(_10697_), .Y(_10715_) );
OAI21X1 OAI21X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_9756_), .B(_9123_), .C(_9759_), .Y(_10716_) );
AOI21X1 AOI21X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_10210_), .B(_10716_), .C(_10209_), .Y(_10717_) );
INVX1 INVX1_1469 ( .gnd(gnd), .vdd(vdd), .A(_10206_), .Y(_10718_) );
INVX1 INVX1_1470 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf2_), .Y(_10720_) );
AOI21X1 AOI21X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_10203_), .B(_10201_), .C(_10198_), .Y(_10721_) );
NOR2X1 NOR2X1_850 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf3_), .B(_10195_), .Y(_10722_) );
INVX1 INVX1_1471 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf0_), .Y(_10723_) );
XNOR2X1 XNOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_12588_), .B(_10636_), .Y(_10724_) );
INVX1 INVX1_1472 ( .gnd(gnd), .vdd(vdd), .A(_10724_), .Y(_10725_) );
OAI21X1 OAI21X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_10189_), .B(_10171_), .C(_10187_), .Y(_10726_) );
XNOR2X1 XNOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_12564_), .B(_10614_), .Y(_10727_) );
INVX1 INVX1_1473 ( .gnd(gnd), .vdd(vdd), .A(_10727_), .Y(_10728_) );
AOI21X1 AOI21X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_9643_), .B(_9101_), .C(_9647_), .Y(_10729_) );
OAI21X1 OAI21X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_10729_), .B(_10181_), .C(_10179_), .Y(_10731_) );
INVX1 INVX1_1474 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_28_), .Y(_10732_) );
XNOR2X1 XNOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_0_), .B(module_2_W_12_), .Y(_10733_) );
XOR2X1 XOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_10733_), .B(module_2_W_8_), .Y(_10734_) );
NAND2X1 NAND2X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_10732_), .B(_10734_), .Y(_10735_) );
XNOR2X1 XNOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_10733_), .B(module_2_W_8_), .Y(_10736_) );
NAND2X1 NAND2X1_1414 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_28_), .B(_10736_), .Y(_10737_) );
NAND3X1 NAND3X1_2379 ( .gnd(gnd), .vdd(vdd), .A(_10175_), .B(_10737_), .C(_10735_), .Y(_10738_) );
AOI21X1 AOI21X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_10737_), .B(_10735_), .C(_10175_), .Y(_10739_) );
INVX2 INVX2_378 ( .gnd(gnd), .vdd(vdd), .A(_10739_), .Y(_10740_) );
AOI21X1 AOI21X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_10738_), .B(_10740_), .C(_10731_), .Y(_10742_) );
INVX1 INVX1_1475 ( .gnd(gnd), .vdd(vdd), .A(_10179_), .Y(_10743_) );
AOI21X1 AOI21X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_10180_), .B(_10174_), .C(_10743_), .Y(_10744_) );
INVX2 INVX2_379 ( .gnd(gnd), .vdd(vdd), .A(_10738_), .Y(_10745_) );
NOR3X1 NOR3X1_307 ( .gnd(gnd), .vdd(vdd), .A(_10744_), .B(_10739_), .C(_10745_), .Y(_10746_) );
OAI21X1 OAI21X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_10746_), .B(_10742_), .C(_10728_), .Y(_10747_) );
OAI21X1 OAI21X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_10745_), .B(_10739_), .C(_10744_), .Y(_10748_) );
NAND3X1 NAND3X1_2380 ( .gnd(gnd), .vdd(vdd), .A(_10731_), .B(_10738_), .C(_10740_), .Y(_10749_) );
NAND3X1 NAND3X1_2381 ( .gnd(gnd), .vdd(vdd), .A(_10727_), .B(_10749_), .C(_10748_), .Y(_10750_) );
NAND3X1 NAND3X1_2382 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf1_), .B(_10750_), .C(_10747_), .Y(_10751_) );
INVX1 INVX1_1476 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf0_), .Y(_10753_) );
NAND3X1 NAND3X1_2383 ( .gnd(gnd), .vdd(vdd), .A(_10728_), .B(_10749_), .C(_10748_), .Y(_10754_) );
OAI21X1 OAI21X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_10746_), .B(_10742_), .C(_10727_), .Y(_10755_) );
NAND3X1 NAND3X1_2384 ( .gnd(gnd), .vdd(vdd), .A(_10753_), .B(_10754_), .C(_10755_), .Y(_10756_) );
NAND3X1 NAND3X1_2385 ( .gnd(gnd), .vdd(vdd), .A(_10183_), .B(_10751_), .C(_10756_), .Y(_10757_) );
INVX1 INVX1_1477 ( .gnd(gnd), .vdd(vdd), .A(_10183_), .Y(_10758_) );
NAND3X1 NAND3X1_2386 ( .gnd(gnd), .vdd(vdd), .A(_10753_), .B(_10750_), .C(_10747_), .Y(_10759_) );
NAND3X1 NAND3X1_2387 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf3_), .B(_10754_), .C(_10755_), .Y(_10760_) );
NAND3X1 NAND3X1_2388 ( .gnd(gnd), .vdd(vdd), .A(_10758_), .B(_10759_), .C(_10760_), .Y(_10761_) );
AOI21X1 AOI21X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_10757_), .B(_10761_), .C(_10726_), .Y(_10762_) );
INVX1 INVX1_1478 ( .gnd(gnd), .vdd(vdd), .A(_10187_), .Y(_10764_) );
AOI21X1 AOI21X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_10188_), .B(_10194_), .C(_10764_), .Y(_10765_) );
AOI21X1 AOI21X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_10759_), .B(_10760_), .C(_10758_), .Y(_10766_) );
AOI21X1 AOI21X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_10751_), .B(_10756_), .C(_10183_), .Y(_10767_) );
NOR3X1 NOR3X1_308 ( .gnd(gnd), .vdd(vdd), .A(_10766_), .B(_10765_), .C(_10767_), .Y(_10768_) );
OAI21X1 OAI21X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_10768_), .B(_10762_), .C(_10725_), .Y(_10769_) );
OAI21X1 OAI21X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_10766_), .B(_10767_), .C(_10765_), .Y(_10770_) );
NAND3X1 NAND3X1_2389 ( .gnd(gnd), .vdd(vdd), .A(_10757_), .B(_10761_), .C(_10726_), .Y(_10771_) );
NAND3X1 NAND3X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_10724_), .B(_10770_), .C(_10771_), .Y(_10772_) );
NAND3X1 NAND3X1_2391 ( .gnd(gnd), .vdd(vdd), .A(_10723_), .B(_10772_), .C(_10769_), .Y(_10773_) );
NAND3X1 NAND3X1_2392 ( .gnd(gnd), .vdd(vdd), .A(_10725_), .B(_10770_), .C(_10771_), .Y(_10775_) );
OAI21X1 OAI21X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_10768_), .B(_10762_), .C(_10724_), .Y(_10776_) );
NAND3X1 NAND3X1_2393 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf4_), .B(_10775_), .C(_10776_), .Y(_10777_) );
AOI21X1 AOI21X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_10773_), .B(_10777_), .C(_10722_), .Y(_10778_) );
INVX1 INVX1_1479 ( .gnd(gnd), .vdd(vdd), .A(_10722_), .Y(_10779_) );
NAND3X1 NAND3X1_2394 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf3_), .B(_10772_), .C(_10769_), .Y(_10780_) );
NAND3X1 NAND3X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_10723_), .B(_10775_), .C(_10776_), .Y(_10781_) );
AOI21X1 AOI21X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_10780_), .B(_10781_), .C(_10779_), .Y(_10782_) );
OAI21X1 OAI21X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_10778_), .B(_10782_), .C(_10721_), .Y(_10783_) );
OAI21X1 OAI21X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_10169_), .B(_10199_), .C(_10202_), .Y(_10784_) );
NAND3X1 NAND3X1_2396 ( .gnd(gnd), .vdd(vdd), .A(_10779_), .B(_10780_), .C(_10781_), .Y(_10786_) );
NAND3X1 NAND3X1_2397 ( .gnd(gnd), .vdd(vdd), .A(_10722_), .B(_10773_), .C(_10777_), .Y(_10787_) );
NAND3X1 NAND3X1_2398 ( .gnd(gnd), .vdd(vdd), .A(_10786_), .B(_10787_), .C(_10784_), .Y(_10788_) );
XNOR2X1 XNOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_10667_), .Y(_10789_) );
NAND3X1 NAND3X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_10789_), .B(_10788_), .C(_10783_), .Y(_10790_) );
AOI21X1 AOI21X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_10786_), .B(_10787_), .C(_10784_), .Y(_10791_) );
NOR3X1 NOR3X1_309 ( .gnd(gnd), .vdd(vdd), .A(_10778_), .B(_10782_), .C(_10721_), .Y(_10792_) );
INVX1 INVX1_1480 ( .gnd(gnd), .vdd(vdd), .A(_10789_), .Y(_10793_) );
OAI21X1 OAI21X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_10792_), .B(_10791_), .C(_10793_), .Y(_10794_) );
NAND3X1 NAND3X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_10720_), .B(_10790_), .C(_10794_), .Y(_10795_) );
NAND3X1 NAND3X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_10793_), .B(_10788_), .C(_10783_), .Y(_10797_) );
OAI21X1 OAI21X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_10792_), .B(_10791_), .C(_10789_), .Y(_10798_) );
NAND3X1 NAND3X1_2402 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf1_), .B(_10797_), .C(_10798_), .Y(_10799_) );
AOI21X1 AOI21X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_10795_), .B(_10799_), .C(_10718_), .Y(_10800_) );
NAND3X1 NAND3X1_2403 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf0_), .B(_10790_), .C(_10794_), .Y(_10801_) );
NAND3X1 NAND3X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_10720_), .B(_10797_), .C(_10798_), .Y(_10802_) );
AOI21X1 AOI21X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_10801_), .B(_10802_), .C(_10206_), .Y(_10803_) );
OAI21X1 OAI21X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_10800_), .B(_10803_), .C(_10717_), .Y(_10804_) );
INVX1 INVX1_1481 ( .gnd(gnd), .vdd(vdd), .A(_10209_), .Y(_10805_) );
OAI21X1 OAI21X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_10166_), .B(_10211_), .C(_10805_), .Y(_10806_) );
NAND3X1 NAND3X1_2405 ( .gnd(gnd), .vdd(vdd), .A(_10206_), .B(_10801_), .C(_10802_), .Y(_10808_) );
NAND3X1 NAND3X1_2406 ( .gnd(gnd), .vdd(vdd), .A(_10718_), .B(_10795_), .C(_10799_), .Y(_10809_) );
NAND3X1 NAND3X1_2407 ( .gnd(gnd), .vdd(vdd), .A(_10808_), .B(_10809_), .C(_10806_), .Y(_10810_) );
NAND3X1 NAND3X1_2408 ( .gnd(gnd), .vdd(vdd), .A(_10715_), .B(_10804_), .C(_10810_), .Y(_10811_) );
INVX1 INVX1_1482 ( .gnd(gnd), .vdd(vdd), .A(_10715_), .Y(_10812_) );
AOI21X1 AOI21X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_10808_), .B(_10809_), .C(_10806_), .Y(_10813_) );
NOR3X1 NOR3X1_310 ( .gnd(gnd), .vdd(vdd), .A(_10800_), .B(_10803_), .C(_10717_), .Y(_10814_) );
OAI21X1 OAI21X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_10814_), .B(_10813_), .C(_10812_), .Y(_10815_) );
NAND3X1 NAND3X1_2409 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf1_), .B(_10811_), .C(_10815_), .Y(_10816_) );
INVX1 INVX1_1483 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf0_), .Y(_10817_) );
NAND3X1 NAND3X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_10812_), .B(_10804_), .C(_10810_), .Y(_10819_) );
OAI21X1 OAI21X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_10814_), .B(_10813_), .C(_10715_), .Y(_10820_) );
NAND3X1 NAND3X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_10817_), .B(_10819_), .C(_10820_), .Y(_10821_) );
NAND3X1 NAND3X1_2412 ( .gnd(gnd), .vdd(vdd), .A(_10221_), .B(_10816_), .C(_10821_), .Y(_10822_) );
INVX1 INVX1_1484 ( .gnd(gnd), .vdd(vdd), .A(_10221_), .Y(_10823_) );
NAND3X1 NAND3X1_2413 ( .gnd(gnd), .vdd(vdd), .A(_10817_), .B(_10811_), .C(_10815_), .Y(_10824_) );
NAND3X1 NAND3X1_2414 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf3_), .B(_10819_), .C(_10820_), .Y(_10825_) );
NAND3X1 NAND3X1_2415 ( .gnd(gnd), .vdd(vdd), .A(_10823_), .B(_10824_), .C(_10825_), .Y(_10826_) );
AOI21X1 AOI21X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_10822_), .B(_10826_), .C(_10714_), .Y(_10827_) );
AOI21X1 AOI21X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_10222_), .B(_10221_), .C(_9796_), .Y(_10828_) );
AOI21X1 AOI21X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_10165_), .B(_10223_), .C(_10828_), .Y(_10830_) );
AOI21X1 AOI21X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_10824_), .B(_10825_), .C(_10823_), .Y(_10831_) );
AOI21X1 AOI21X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_10816_), .B(_10821_), .C(_10221_), .Y(_10832_) );
NOR3X1 NOR3X1_311 ( .gnd(gnd), .vdd(vdd), .A(_10831_), .B(_10832_), .C(_10830_), .Y(_10833_) );
OAI21X1 OAI21X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_10833_), .B(_10827_), .C(_10711_), .Y(_10834_) );
INVX1 INVX1_1485 ( .gnd(gnd), .vdd(vdd), .A(_10711_), .Y(_10835_) );
OAI21X1 OAI21X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_10831_), .B(_10832_), .C(_10830_), .Y(_10836_) );
NAND3X1 NAND3X1_2416 ( .gnd(gnd), .vdd(vdd), .A(_10822_), .B(_10826_), .C(_10714_), .Y(_10837_) );
NAND3X1 NAND3X1_2417 ( .gnd(gnd), .vdd(vdd), .A(_10835_), .B(_10836_), .C(_10837_), .Y(_10838_) );
NAND3X1 NAND3X1_2418 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf2_), .B(_10838_), .C(_10834_), .Y(_10839_) );
INVX1 INVX1_1486 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf1_), .Y(_10841_) );
NAND3X1 NAND3X1_2419 ( .gnd(gnd), .vdd(vdd), .A(_10711_), .B(_10836_), .C(_10837_), .Y(_10842_) );
OAI21X1 OAI21X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_10833_), .B(_10827_), .C(_10835_), .Y(_10843_) );
NAND3X1 NAND3X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_10841_), .B(_10842_), .C(_10843_), .Y(_10844_) );
NAND3X1 NAND3X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_10232_), .B(_10839_), .C(_10844_), .Y(_10845_) );
INVX1 INVX1_1487 ( .gnd(gnd), .vdd(vdd), .A(_10232_), .Y(_10846_) );
NAND3X1 NAND3X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_10841_), .B(_10838_), .C(_10834_), .Y(_10847_) );
NAND3X1 NAND3X1_2423 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf0_), .B(_10842_), .C(_10843_), .Y(_10848_) );
NAND3X1 NAND3X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_10846_), .B(_10847_), .C(_10848_), .Y(_10849_) );
AOI21X1 AOI21X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_10845_), .B(_10849_), .C(_10710_), .Y(_10850_) );
INVX1 INVX1_1488 ( .gnd(gnd), .vdd(vdd), .A(_10231_), .Y(_10852_) );
AOI21X1 AOI21X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_10234_), .B(_10163_), .C(_10852_), .Y(_10853_) );
AOI21X1 AOI21X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_10847_), .B(_10848_), .C(_10846_), .Y(_10854_) );
AOI21X1 AOI21X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_10839_), .B(_10844_), .C(_10232_), .Y(_10855_) );
NOR3X1 NOR3X1_312 ( .gnd(gnd), .vdd(vdd), .A(_10854_), .B(_10853_), .C(_10855_), .Y(_10856_) );
OAI21X1 OAI21X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_10856_), .B(_10850_), .C(_10709_), .Y(_10857_) );
INVX1 INVX1_1489 ( .gnd(gnd), .vdd(vdd), .A(_10709_), .Y(_10858_) );
OAI21X1 OAI21X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_10854_), .B(_10855_), .C(_10853_), .Y(_10859_) );
NAND3X1 NAND3X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_10845_), .B(_10849_), .C(_10710_), .Y(_10860_) );
NAND3X1 NAND3X1_2426 ( .gnd(gnd), .vdd(vdd), .A(_10858_), .B(_10860_), .C(_10859_), .Y(_10861_) );
NAND3X1 NAND3X1_2427 ( .gnd(gnd), .vdd(vdd), .A(_10707_), .B(_10861_), .C(_10857_), .Y(_10863_) );
NAND3X1 NAND3X1_2428 ( .gnd(gnd), .vdd(vdd), .A(_10709_), .B(_10860_), .C(_10859_), .Y(_10864_) );
OAI21X1 OAI21X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_10856_), .B(_10850_), .C(_10858_), .Y(_10865_) );
NAND3X1 NAND3X1_2429 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf2_), .B(_10864_), .C(_10865_), .Y(_10866_) );
AOI21X1 AOI21X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_10863_), .B(_10866_), .C(_10706_), .Y(_10867_) );
NAND3X1 NAND3X1_2430 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf1_), .B(_10861_), .C(_10857_), .Y(_10868_) );
NAND3X1 NAND3X1_2431 ( .gnd(gnd), .vdd(vdd), .A(_10707_), .B(_10864_), .C(_10865_), .Y(_10869_) );
AOI21X1 AOI21X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_10868_), .B(_10869_), .C(_10243_), .Y(_10870_) );
OAI21X1 OAI21X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_10867_), .B(_10870_), .C(_10705_), .Y(_10871_) );
NAND2X1 NAND2X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_10242_), .B(_10246_), .Y(_10872_) );
NAND3X1 NAND3X1_2432 ( .gnd(gnd), .vdd(vdd), .A(_10243_), .B(_10868_), .C(_10869_), .Y(_10874_) );
NAND3X1 NAND3X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_10706_), .B(_10863_), .C(_10866_), .Y(_10875_) );
NAND3X1 NAND3X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_10872_), .B(_10874_), .C(_10875_), .Y(_10876_) );
NAND3X1 NAND3X1_2435 ( .gnd(gnd), .vdd(vdd), .A(_11180_), .B(_10876_), .C(_10871_), .Y(_10877_) );
AOI21X1 AOI21X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_10874_), .B(_10875_), .C(_10872_), .Y(_10878_) );
NOR3X1 NOR3X1_313 ( .gnd(gnd), .vdd(vdd), .A(_10870_), .B(_10705_), .C(_10867_), .Y(_10879_) );
OAI21X1 OAI21X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_10879_), .B(_10878_), .C(_10796_), .Y(_10880_) );
NAND2X1 NAND2X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_10877_), .B(_10880_), .Y(_10881_) );
NAND3X1 NAND3X1_2436 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_140_), .B(_8902_), .C(_10881_), .Y(_10882_) );
INVX1 INVX1_1490 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_140_), .Y(_10883_) );
OAI21X1 OAI21X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_10879_), .B(_10878_), .C(_11180_), .Y(_10885_) );
NAND3X1 NAND3X1_2437 ( .gnd(gnd), .vdd(vdd), .A(_10796_), .B(_10876_), .C(_10871_), .Y(_10886_) );
NAND3X1 NAND3X1_2438 ( .gnd(gnd), .vdd(vdd), .A(_8902_), .B(_10886_), .C(_10885_), .Y(_10887_) );
NAND2X1 NAND2X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_10883_), .B(_10887_), .Y(_10888_) );
AOI21X1 AOI21X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_10882_), .B(_10888_), .C(_10704_), .Y(_10889_) );
INVX1 INVX1_1491 ( .gnd(gnd), .vdd(vdd), .A(_10704_), .Y(_10890_) );
NAND2X1 NAND2X1_1418 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_140_), .B(_10887_), .Y(_10891_) );
NAND3X1 NAND3X1_2439 ( .gnd(gnd), .vdd(vdd), .A(_10883_), .B(_8902_), .C(_10881_), .Y(_10892_) );
AOI21X1 AOI21X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_10891_), .B(_10892_), .C(_10890_), .Y(_10893_) );
OAI21X1 OAI21X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_10893_), .B(_10889_), .C(_10703_), .Y(_10894_) );
NAND3X1 NAND3X1_2440 ( .gnd(gnd), .vdd(vdd), .A(_10890_), .B(_10891_), .C(_10892_), .Y(_10896_) );
NAND3X1 NAND3X1_2441 ( .gnd(gnd), .vdd(vdd), .A(_10704_), .B(_10882_), .C(_10888_), .Y(_10897_) );
NAND3X1 NAND3X1_2442 ( .gnd(gnd), .vdd(vdd), .A(_10702_), .B(_10896_), .C(_10897_), .Y(_10898_) );
NAND3X1 NAND3X1_2443 ( .gnd(gnd), .vdd(vdd), .A(_10829_), .B(_10898_), .C(_10894_), .Y(_10899_) );
NAND2X1 NAND2X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_10898_), .B(_10894_), .Y(_10900_) );
AOI21X1 AOI21X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_11147_), .B(_10900_), .C(_8931_), .Y(_10901_) );
NAND3X1 NAND3X1_2444 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_156_), .B(_10899_), .C(_10901_), .Y(_10902_) );
INVX1 INVX1_1492 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_156_), .Y(_10903_) );
AOI21X1 AOI21X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_10896_), .B(_10897_), .C(_10702_), .Y(_10904_) );
NOR3X1 NOR3X1_314 ( .gnd(gnd), .vdd(vdd), .A(_10889_), .B(_10893_), .C(_10703_), .Y(_10905_) );
OAI21X1 OAI21X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_10905_), .B(_10904_), .C(_11147_), .Y(_10907_) );
NAND3X1 NAND3X1_2445 ( .gnd(gnd), .vdd(vdd), .A(_8928_), .B(_10899_), .C(_10907_), .Y(_10908_) );
NAND2X1 NAND2X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_10903_), .B(_10908_), .Y(_10909_) );
AOI21X1 AOI21X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_10902_), .B(_10909_), .C(_10263_), .Y(_10910_) );
NAND2X1 NAND2X1_1421 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_156_), .B(_10908_), .Y(_10911_) );
NAND3X1 NAND3X1_2446 ( .gnd(gnd), .vdd(vdd), .A(_10903_), .B(_10899_), .C(_10901_), .Y(_10912_) );
AOI21X1 AOI21X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_10912_), .B(_10911_), .C(_10261_), .Y(_10913_) );
OAI21X1 OAI21X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_10913_), .B(_10910_), .C(_10701_), .Y(_10914_) );
NAND3X1 NAND3X1_2447 ( .gnd(gnd), .vdd(vdd), .A(_9945_), .B(_10259_), .C(_10263_), .Y(_10915_) );
OAI21X1 OAI21X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_10267_), .B(_10264_), .C(_10915_), .Y(_10916_) );
NAND3X1 NAND3X1_2448 ( .gnd(gnd), .vdd(vdd), .A(_10261_), .B(_10912_), .C(_10911_), .Y(_10918_) );
NAND3X1 NAND3X1_2449 ( .gnd(gnd), .vdd(vdd), .A(_10263_), .B(_10902_), .C(_10909_), .Y(_10919_) );
NAND3X1 NAND3X1_2450 ( .gnd(gnd), .vdd(vdd), .A(_10916_), .B(_10918_), .C(_10919_), .Y(_10920_) );
AOI21X1 AOI21X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_10920_), .B(_10914_), .C(_10862_), .Y(_10921_) );
NAND2X1 NAND2X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_10920_), .B(_10914_), .Y(_10922_) );
OAI21X1 OAI21X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_10922_), .B(_11114_), .C(_8953_), .Y(_10923_) );
OAI21X1 OAI21X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_10923_), .B(_10921_), .C(module_2_W_172_), .Y(_10924_) );
INVX1 INVX1_1493 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_172_), .Y(_10925_) );
NAND3X1 NAND3X1_2451 ( .gnd(gnd), .vdd(vdd), .A(_11114_), .B(_10920_), .C(_10914_), .Y(_10926_) );
AOI21X1 AOI21X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_10918_), .B(_10919_), .C(_10916_), .Y(_10927_) );
NOR3X1 NOR3X1_315 ( .gnd(gnd), .vdd(vdd), .A(_10910_), .B(_10701_), .C(_10913_), .Y(_10929_) );
OAI21X1 OAI21X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_10929_), .B(_10927_), .C(_10862_), .Y(_10930_) );
NAND2X1 NAND2X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_10926_), .B(_10930_), .Y(_10931_) );
NAND3X1 NAND3X1_2452 ( .gnd(gnd), .vdd(vdd), .A(_10925_), .B(_8953_), .C(_10931_), .Y(_10932_) );
NAND3X1 NAND3X1_2453 ( .gnd(gnd), .vdd(vdd), .A(_10699_), .B(_10924_), .C(_10932_), .Y(_10933_) );
NAND3X1 NAND3X1_2454 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_172_), .B(_8953_), .C(_10931_), .Y(_10934_) );
OAI21X1 OAI21X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_10923_), .B(_10921_), .C(_10925_), .Y(_10935_) );
NAND3X1 NAND3X1_2455 ( .gnd(gnd), .vdd(vdd), .A(_10272_), .B(_10935_), .C(_10934_), .Y(_10936_) );
AOI21X1 AOI21X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_10933_), .B(_10936_), .C(_10698_), .Y(_10937_) );
INVX1 INVX1_1494 ( .gnd(gnd), .vdd(vdd), .A(_10275_), .Y(_10938_) );
AOI21X1 AOI21X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_10938_), .B(_10155_), .C(_10274_), .Y(_10940_) );
AOI21X1 AOI21X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_10935_), .B(_10934_), .C(_10272_), .Y(_10941_) );
AOI21X1 AOI21X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_10924_), .B(_10932_), .C(_10699_), .Y(_10942_) );
NOR3X1 NOR3X1_316 ( .gnd(gnd), .vdd(vdd), .A(_10941_), .B(_10942_), .C(_10940_), .Y(_10943_) );
OAI21X1 OAI21X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_10943_), .B(_10937_), .C(_11092_), .Y(_10944_) );
OAI21X1 OAI21X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_10942_), .B(_10941_), .C(_10940_), .Y(_10945_) );
NAND3X1 NAND3X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_10698_), .B(_10933_), .C(_10936_), .Y(_10946_) );
NAND3X1 NAND3X1_2457 ( .gnd(gnd), .vdd(vdd), .A(_10895_), .B(_10946_), .C(_10945_), .Y(_10947_) );
NAND3X1 NAND3X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_8972_), .B(_10947_), .C(_10944_), .Y(_10948_) );
NAND2X1 NAND2X1_1424 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_188_), .B(_10948_), .Y(_10949_) );
INVX1 INVX1_1495 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_188_), .Y(_10951_) );
NAND3X1 NAND3X1_2459 ( .gnd(gnd), .vdd(vdd), .A(_11092_), .B(_10946_), .C(_10945_), .Y(_10952_) );
OAI21X1 OAI21X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_10943_), .B(_10937_), .C(_10895_), .Y(_10953_) );
NAND2X1 NAND2X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_10952_), .B(_10953_), .Y(_10954_) );
NAND3X1 NAND3X1_2460 ( .gnd(gnd), .vdd(vdd), .A(_10951_), .B(_8972_), .C(_10954_), .Y(_10955_) );
NAND3X1 NAND3X1_2461 ( .gnd(gnd), .vdd(vdd), .A(_10695_), .B(_10949_), .C(_10955_), .Y(_10956_) );
NAND3X1 NAND3X1_2462 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_188_), .B(_8972_), .C(_10954_), .Y(_10957_) );
NAND2X1 NAND2X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_10951_), .B(_10948_), .Y(_10958_) );
NAND3X1 NAND3X1_2463 ( .gnd(gnd), .vdd(vdd), .A(_10282_), .B(_10957_), .C(_10958_), .Y(_10959_) );
AOI21X1 AOI21X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_10956_), .B(_10959_), .C(_10694_), .Y(_10960_) );
INVX1 INVX1_1496 ( .gnd(gnd), .vdd(vdd), .A(_10285_), .Y(_10962_) );
AOI21X1 AOI21X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_10152_), .B(_10962_), .C(_10284_), .Y(_10963_) );
AOI21X1 AOI21X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_10957_), .B(_10958_), .C(_10282_), .Y(_10964_) );
AOI21X1 AOI21X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_10949_), .B(_10955_), .C(_10695_), .Y(_10965_) );
NOR3X1 NOR3X1_317 ( .gnd(gnd), .vdd(vdd), .A(_10964_), .B(_10965_), .C(_10963_), .Y(_10966_) );
OAI21X1 OAI21X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_10966_), .B(_10960_), .C(_10928_), .Y(_10967_) );
OAI21X1 OAI21X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_10965_), .B(_10964_), .C(_10963_), .Y(_10968_) );
NAND3X1 NAND3X1_2464 ( .gnd(gnd), .vdd(vdd), .A(_10694_), .B(_10956_), .C(_10959_), .Y(_10969_) );
NAND3X1 NAND3X1_2465 ( .gnd(gnd), .vdd(vdd), .A(_11059_), .B(_10969_), .C(_10968_), .Y(_10970_) );
NAND2X1 NAND2X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_10970_), .B(_10967_), .Y(_10971_) );
NAND3X1 NAND3X1_2466 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_204_), .B(_8999_), .C(_10971_), .Y(_10973_) );
INVX1 INVX1_1497 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_204_), .Y(_10974_) );
AOI21X1 AOI21X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_10969_), .B(_10968_), .C(_10928_), .Y(_10975_) );
NAND2X1 NAND2X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_10969_), .B(_10968_), .Y(_10976_) );
OAI21X1 OAI21X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_10976_), .B(_11059_), .C(_8999_), .Y(_10977_) );
OAI21X1 OAI21X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_10977_), .B(_10975_), .C(_10974_), .Y(_10978_) );
AOI21X1 AOI21X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_10978_), .B(_10973_), .C(_10293_), .Y(_10979_) );
OAI21X1 OAI21X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_10977_), .B(_10975_), .C(module_2_W_204_), .Y(_10980_) );
NAND3X1 NAND3X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_10974_), .B(_8999_), .C(_10971_), .Y(_10981_) );
AOI21X1 AOI21X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_10980_), .B(_10981_), .C(_10292_), .Y(_10982_) );
OAI21X1 OAI21X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_10982_), .B(_10979_), .C(_10693_), .Y(_10984_) );
AOI21X1 AOI21X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_10291_), .B(_10293_), .C(_10055_), .Y(_10985_) );
OAI21X1 OAI21X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_10985_), .B(_10150_), .C(_10294_), .Y(_10986_) );
NAND3X1 NAND3X1_2468 ( .gnd(gnd), .vdd(vdd), .A(_10292_), .B(_10980_), .C(_10981_), .Y(_10987_) );
NAND3X1 NAND3X1_2469 ( .gnd(gnd), .vdd(vdd), .A(_10293_), .B(_10978_), .C(_10973_), .Y(_10988_) );
NAND3X1 NAND3X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_10987_), .B(_10988_), .C(_10986_), .Y(_10989_) );
NAND3X1 NAND3X1_2471 ( .gnd(gnd), .vdd(vdd), .A(_11038_), .B(_10989_), .C(_10984_), .Y(_10990_) );
AOI21X1 AOI21X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_10987_), .B(_10988_), .C(_10986_), .Y(_10991_) );
NOR3X1 NOR3X1_318 ( .gnd(gnd), .vdd(vdd), .A(_10979_), .B(_10693_), .C(_10982_), .Y(_10992_) );
OAI21X1 OAI21X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_10992_), .B(_10991_), .C(_10961_), .Y(_10993_) );
NAND2X1 NAND2X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_10990_), .B(_10993_), .Y(_10995_) );
NAND3X1 NAND3X1_2472 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_220_), .B(_9020_), .C(_10995_), .Y(_10996_) );
INVX1 INVX1_1498 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_220_), .Y(_10997_) );
AOI21X1 AOI21X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_10989_), .B(_10984_), .C(_10961_), .Y(_10998_) );
NAND2X1 NAND2X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_10989_), .B(_10984_), .Y(_10999_) );
OAI21X1 OAI21X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_10999_), .B(_11038_), .C(_9020_), .Y(_11000_) );
OAI21X1 OAI21X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_11000_), .B(_10998_), .C(_10997_), .Y(_11001_) );
AOI21X1 AOI21X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_11001_), .B(_10996_), .C(_10306_), .Y(_11002_) );
OAI21X1 OAI21X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_11000_), .B(_10998_), .C(module_2_W_220_), .Y(_11003_) );
NAND3X1 NAND3X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_10997_), .B(_9020_), .C(_10995_), .Y(_11004_) );
AOI21X1 AOI21X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_11003_), .B(_11004_), .C(_10303_), .Y(_11006_) );
OAI21X1 OAI21X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_11002_), .B(_11006_), .C(_10691_), .Y(_11007_) );
AOI21X1 AOI21X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_10089_), .B(_10097_), .C(_10099_), .Y(_11008_) );
NAND3X1 NAND3X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_10092_), .B(_10306_), .C(_10305_), .Y(_11009_) );
OAI21X1 OAI21X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_11008_), .B(_10307_), .C(_11009_), .Y(_11010_) );
NAND3X1 NAND3X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_10303_), .B(_11003_), .C(_11004_), .Y(_11011_) );
NAND3X1 NAND3X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_10306_), .B(_11001_), .C(_10996_), .Y(_11012_) );
NAND3X1 NAND3X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_11010_), .B(_11011_), .C(_11012_), .Y(_11013_) );
AOI21X1 AOI21X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_11013_), .B(_11007_), .C(_10994_), .Y(_11014_) );
NAND2X1 NAND2X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_11013_), .B(_11007_), .Y(_11015_) );
OAI21X1 OAI21X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_11015_), .B(_11005_), .C(_9046_), .Y(_11017_) );
OAI21X1 OAI21X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_11017_), .B(_11014_), .C(module_2_W_236_), .Y(_11018_) );
INVX1 INVX1_1499 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_236_), .Y(_11019_) );
NAND3X1 NAND3X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_11005_), .B(_11013_), .C(_11007_), .Y(_11020_) );
AOI21X1 AOI21X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_11011_), .B(_11012_), .C(_11010_), .Y(_11021_) );
NOR3X1 NOR3X1_319 ( .gnd(gnd), .vdd(vdd), .A(_11002_), .B(_10691_), .C(_11006_), .Y(_11022_) );
OAI21X1 OAI21X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_11022_), .B(_11021_), .C(_10994_), .Y(_11023_) );
NAND2X1 NAND2X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_11020_), .B(_11023_), .Y(_11024_) );
NAND3X1 NAND3X1_2479 ( .gnd(gnd), .vdd(vdd), .A(_11019_), .B(_9046_), .C(_11024_), .Y(_11025_) );
NAND3X1 NAND3X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_10689_), .B(_11018_), .C(_11025_), .Y(_11026_) );
NAND3X1 NAND3X1_2481 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_236_), .B(_9046_), .C(_11024_), .Y(_11028_) );
OAI21X1 OAI21X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_11017_), .B(_11014_), .C(_11019_), .Y(_11029_) );
NAND3X1 NAND3X1_2482 ( .gnd(gnd), .vdd(vdd), .A(_10313_), .B(_11029_), .C(_11028_), .Y(_11030_) );
AOI21X1 AOI21X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_11026_), .B(_11030_), .C(_10688_), .Y(_11031_) );
INVX1 INVX1_1500 ( .gnd(gnd), .vdd(vdd), .A(_10316_), .Y(_11032_) );
AOI21X1 AOI21X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_10319_), .B(_11032_), .C(_10315_), .Y(_11033_) );
NAND3X1 NAND3X1_2483 ( .gnd(gnd), .vdd(vdd), .A(_10689_), .B(_11029_), .C(_11028_), .Y(_11034_) );
NAND3X1 NAND3X1_2484 ( .gnd(gnd), .vdd(vdd), .A(_10313_), .B(_11018_), .C(_11025_), .Y(_11035_) );
AOI21X1 AOI21X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_11034_), .B(_11035_), .C(_11033_), .Y(_11036_) );
OAI21X1 OAI21X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_11036_), .B(_11031_), .C(_12239_), .Y(_11037_) );
AOI21X1 AOI21X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_11029_), .B(_11028_), .C(_10313_), .Y(_11039_) );
AOI21X1 AOI21X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_11018_), .B(_11025_), .C(_10689_), .Y(_11040_) );
OAI21X1 OAI21X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_11039_), .B(_11040_), .C(_11033_), .Y(_11041_) );
NAND3X1 NAND3X1_2485 ( .gnd(gnd), .vdd(vdd), .A(_10688_), .B(_11026_), .C(_11030_), .Y(_11042_) );
NAND3X1 NAND3X1_2486 ( .gnd(gnd), .vdd(vdd), .A(_12240_), .B(_11042_), .C(_11041_), .Y(_11043_) );
NAND2X1 NAND2X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_11043_), .B(_11037_), .Y(_11044_) );
NAND3X1 NAND3X1_2487 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_252_), .B(_9070_), .C(_11044_), .Y(_11045_) );
INVX1 INVX1_1501 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_252_), .Y(_11046_) );
AOI21X1 AOI21X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_11042_), .B(_11041_), .C(_12239_), .Y(_11047_) );
NAND2X1 NAND2X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_11042_), .B(_11041_), .Y(_11048_) );
OAI21X1 OAI21X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_11048_), .B(_12240_), .C(_9070_), .Y(_11050_) );
OAI21X1 OAI21X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_11050_), .B(_11047_), .C(_11046_), .Y(_11051_) );
AOI21X1 AOI21X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_11051_), .B(_11045_), .C(_10680_), .Y(_11052_) );
INVX1 INVX1_1502 ( .gnd(gnd), .vdd(vdd), .A(_11052_), .Y(_11053_) );
NAND3X1 NAND3X1_2488 ( .gnd(gnd), .vdd(vdd), .A(_10680_), .B(_11051_), .C(_11045_), .Y(_11054_) );
NAND2X1 NAND2X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_11054_), .B(_11053_), .Y(_11055_) );
XOR2X1 XOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_11055_), .B(_10687_), .Y(module_2_H_20_) );
OAI21X1 OAI21X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_11052_), .B(_10687_), .C(_11054_), .Y(_11056_) );
NAND2X1 NAND2X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_9070_), .B(_11044_), .Y(_11057_) );
NOR2X1 NOR2X1_851 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_252_), .B(_11057_), .Y(_11058_) );
AOI21X1 AOI21X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_10688_), .B(_11030_), .C(_11039_), .Y(_11060_) );
INVX1 INVX1_1503 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_237_), .Y(_11061_) );
OAI21X1 OAI21X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_11006_), .B(_10691_), .C(_11011_), .Y(_11062_) );
INVX1 INVX1_1504 ( .gnd(gnd), .vdd(vdd), .A(_11003_), .Y(_11063_) );
AOI21X1 AOI21X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_10988_), .B(_10986_), .C(_10979_), .Y(_11064_) );
INVX1 INVX1_1505 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_205_), .Y(_11065_) );
OAI21X1 OAI21X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_10963_), .B(_10965_), .C(_10956_), .Y(_11066_) );
INVX1 INVX1_1506 ( .gnd(gnd), .vdd(vdd), .A(_10949_), .Y(_11067_) );
AOI21X1 AOI21X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_10698_), .B(_10936_), .C(_10941_), .Y(_11068_) );
INVX1 INVX1_1507 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_173_), .Y(_11069_) );
INVX1 INVX1_1508 ( .gnd(gnd), .vdd(vdd), .A(_12010_), .Y(_11071_) );
AOI21X1 AOI21X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_10916_), .B(_10919_), .C(_10910_), .Y(_11072_) );
INVX1 INVX1_1509 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_157_), .Y(_11073_) );
INVX1 INVX1_1510 ( .gnd(gnd), .vdd(vdd), .A(_11926_), .Y(_11074_) );
AOI21X1 AOI21X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_10702_), .B(_10897_), .C(_10889_), .Y(_11075_) );
INVX1 INVX1_1511 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_141_), .Y(_11076_) );
OAI21X1 OAI21X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_10870_), .B(_10705_), .C(_10874_), .Y(_11077_) );
INVX1 INVX1_1512 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf3_), .Y(_11078_) );
AOI21X1 AOI21X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_10849_), .B(_10710_), .C(_10854_), .Y(_11079_) );
INVX1 INVX1_1513 ( .gnd(gnd), .vdd(vdd), .A(_10847_), .Y(_11080_) );
INVX1 INVX1_1514 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf2_), .Y(_11082_) );
AOI21X1 AOI21X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_10826_), .B(_10714_), .C(_10831_), .Y(_11083_) );
INVX1 INVX1_1515 ( .gnd(gnd), .vdd(vdd), .A(_10824_), .Y(_11084_) );
INVX1 INVX1_1516 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf2_), .Y(_11085_) );
AOI21X1 AOI21X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_10809_), .B(_10806_), .C(_10800_), .Y(_11086_) );
INVX1 INVX1_1517 ( .gnd(gnd), .vdd(vdd), .A(_10795_), .Y(_11087_) );
INVX1 INVX1_1518 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf2_), .Y(_11088_) );
OAI21X1 OAI21X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_10721_), .B(_10782_), .C(_10786_), .Y(_11089_) );
INVX1 INVX1_1519 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf0_), .Y(_11090_) );
AOI21X1 AOI21X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_10761_), .B(_10726_), .C(_10766_), .Y(_11091_) );
INVX1 INVX1_1520 ( .gnd(gnd), .vdd(vdd), .A(_10759_), .Y(_11093_) );
INVX1 INVX1_1521 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf3_), .Y(_11094_) );
OAI21X1 OAI21X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_10745_), .B(_10744_), .C(_10740_), .Y(_11095_) );
INVX1 INVX1_1522 ( .gnd(gnd), .vdd(vdd), .A(_10735_), .Y(_11096_) );
XOR2X1 XOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_12_), .B(module_2_W_13_), .Y(_11097_) );
INVX1 INVX1_1523 ( .gnd(gnd), .vdd(vdd), .A(_11097_), .Y(_11098_) );
OAI21X1 OAI21X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_11378_), .B(_11389_), .C(module_2_W_9_), .Y(_11099_) );
NAND2X1 NAND2X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_9096_), .B(_9239_), .Y(_11100_) );
NAND2X1 NAND2X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_11099_), .B(_11100_), .Y(_11101_) );
NAND2X1 NAND2X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_11098_), .B(_11101_), .Y(_11102_) );
NAND3X1 NAND3X1_2489 ( .gnd(gnd), .vdd(vdd), .A(_11097_), .B(_11099_), .C(_11100_), .Y(_11104_) );
AOI21X1 AOI21X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_11104_), .B(_11102_), .C(module_2_W_29_), .Y(_11105_) );
INVX1 INVX1_1524 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_29_), .Y(_11106_) );
NAND2X1 NAND2X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_11097_), .B(_11101_), .Y(_11107_) );
NAND3X1 NAND3X1_2490 ( .gnd(gnd), .vdd(vdd), .A(_11098_), .B(_11099_), .C(_11100_), .Y(_11108_) );
AOI21X1 AOI21X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_11108_), .B(_11107_), .C(_11106_), .Y(_11109_) );
OAI21X1 OAI21X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_11109_), .B(_11105_), .C(_11096_), .Y(_11110_) );
NAND3X1 NAND3X1_2491 ( .gnd(gnd), .vdd(vdd), .A(_11106_), .B(_11108_), .C(_11107_), .Y(_11111_) );
NAND3X1 NAND3X1_2492 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_29_), .B(_11104_), .C(_11102_), .Y(_11112_) );
NAND3X1 NAND3X1_2493 ( .gnd(gnd), .vdd(vdd), .A(_10735_), .B(_11112_), .C(_11111_), .Y(_11113_) );
NAND3X1 NAND3X1_2494 ( .gnd(gnd), .vdd(vdd), .A(_11110_), .B(_11113_), .C(_11095_), .Y(_11115_) );
AOI21X1 AOI21X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_10738_), .B(_10731_), .C(_10739_), .Y(_11116_) );
AOI21X1 AOI21X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_11112_), .B(_11111_), .C(_10735_), .Y(_11117_) );
NOR3X1 NOR3X1_320 ( .gnd(gnd), .vdd(vdd), .A(_11105_), .B(_11096_), .C(_11109_), .Y(_11118_) );
OAI21X1 OAI21X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_11118_), .B(_11117_), .C(_11116_), .Y(_11119_) );
XNOR2X1 XNOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_9102_), .B(_11465_), .Y(_11120_) );
INVX1 INVX1_1525 ( .gnd(gnd), .vdd(vdd), .A(_11120_), .Y(_11121_) );
NAND3X1 NAND3X1_2495 ( .gnd(gnd), .vdd(vdd), .A(_11119_), .B(_11121_), .C(_11115_), .Y(_11122_) );
NOR3X1 NOR3X1_321 ( .gnd(gnd), .vdd(vdd), .A(_11116_), .B(_11117_), .C(_11118_), .Y(_11123_) );
AOI21X1 AOI21X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_11110_), .B(_11113_), .C(_11095_), .Y(_11124_) );
OAI21X1 OAI21X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_11123_), .B(_11124_), .C(_11120_), .Y(_11126_) );
NAND3X1 NAND3X1_2496 ( .gnd(gnd), .vdd(vdd), .A(_11094_), .B(_11122_), .C(_11126_), .Y(_11127_) );
NAND3X1 NAND3X1_2497 ( .gnd(gnd), .vdd(vdd), .A(_11119_), .B(_11120_), .C(_11115_), .Y(_11128_) );
OAI21X1 OAI21X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_11123_), .B(_11124_), .C(_11121_), .Y(_11129_) );
NAND3X1 NAND3X1_2498 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf2_), .B(_11128_), .C(_11129_), .Y(_11130_) );
NAND3X1 NAND3X1_2499 ( .gnd(gnd), .vdd(vdd), .A(_11093_), .B(_11127_), .C(_11130_), .Y(_11131_) );
AOI21X1 AOI21X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_11128_), .B(_11129_), .C(bloque_datos_13_bF_buf1_), .Y(_11132_) );
AOI21X1 AOI21X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_11122_), .B(_11126_), .C(_11094_), .Y(_11133_) );
OAI21X1 OAI21X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_11132_), .B(_11133_), .C(_10759_), .Y(_11134_) );
NAND3X1 NAND3X1_2500 ( .gnd(gnd), .vdd(vdd), .A(_11131_), .B(_11134_), .C(_11091_), .Y(_11135_) );
OAI21X1 OAI21X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_10767_), .B(_10765_), .C(_10757_), .Y(_11137_) );
NAND3X1 NAND3X1_2501 ( .gnd(gnd), .vdd(vdd), .A(_10759_), .B(_11127_), .C(_11130_), .Y(_11138_) );
OAI21X1 OAI21X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_11132_), .B(_11133_), .C(_11093_), .Y(_11139_) );
NAND3X1 NAND3X1_2502 ( .gnd(gnd), .vdd(vdd), .A(_11138_), .B(_11139_), .C(_11137_), .Y(_11140_) );
XNOR2X1 XNOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_9302_), .B(_11509_), .Y(_11141_) );
INVX1 INVX1_1526 ( .gnd(gnd), .vdd(vdd), .A(_11141_), .Y(_11142_) );
NAND3X1 NAND3X1_2503 ( .gnd(gnd), .vdd(vdd), .A(_11140_), .B(_11142_), .C(_11135_), .Y(_11143_) );
AOI21X1 AOI21X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_11138_), .B(_11139_), .C(_11137_), .Y(_11144_) );
AOI21X1 AOI21X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_11131_), .B(_11134_), .C(_11091_), .Y(_11145_) );
OAI21X1 OAI21X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_11145_), .B(_11144_), .C(_11141_), .Y(_11146_) );
NAND3X1 NAND3X1_2504 ( .gnd(gnd), .vdd(vdd), .A(_11090_), .B(_11143_), .C(_11146_), .Y(_11148_) );
NOR3X1 NOR3X1_322 ( .gnd(gnd), .vdd(vdd), .A(_11144_), .B(_11141_), .C(_11145_), .Y(_11149_) );
AOI21X1 AOI21X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_11140_), .B(_11135_), .C(_11142_), .Y(_11150_) );
OAI21X1 OAI21X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_11149_), .B(_11150_), .C(bloque_datos_29_bF_buf4_), .Y(_11151_) );
NAND3X1 NAND3X1_2505 ( .gnd(gnd), .vdd(vdd), .A(_10773_), .B(_11148_), .C(_11151_), .Y(_11152_) );
INVX1 INVX1_1527 ( .gnd(gnd), .vdd(vdd), .A(_10773_), .Y(_11153_) );
NOR3X1 NOR3X1_323 ( .gnd(gnd), .vdd(vdd), .A(_11150_), .B(bloque_datos_29_bF_buf3_), .C(_11149_), .Y(_11154_) );
AOI21X1 AOI21X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_11143_), .B(_11146_), .C(_11090_), .Y(_11155_) );
OAI21X1 OAI21X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_11154_), .B(_11155_), .C(_11153_), .Y(_11156_) );
AOI21X1 AOI21X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_11152_), .B(_11156_), .C(_11089_), .Y(_11157_) );
AOI21X1 AOI21X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_10787_), .B(_10784_), .C(_10778_), .Y(_11159_) );
NAND3X1 NAND3X1_2506 ( .gnd(gnd), .vdd(vdd), .A(_11153_), .B(_11148_), .C(_11151_), .Y(_11160_) );
OAI21X1 OAI21X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_11154_), .B(_11155_), .C(_10773_), .Y(_11161_) );
AOI21X1 AOI21X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_11160_), .B(_11161_), .C(_11159_), .Y(_11162_) );
XNOR2X1 XNOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_9119_), .B(_11564_), .Y(_11163_) );
NOR3X1 NOR3X1_324 ( .gnd(gnd), .vdd(vdd), .A(_11162_), .B(_11163_), .C(_11157_), .Y(_11164_) );
NAND3X1 NAND3X1_2507 ( .gnd(gnd), .vdd(vdd), .A(_11160_), .B(_11159_), .C(_11161_), .Y(_11165_) );
NAND3X1 NAND3X1_2508 ( .gnd(gnd), .vdd(vdd), .A(_11089_), .B(_11152_), .C(_11156_), .Y(_11166_) );
INVX1 INVX1_1528 ( .gnd(gnd), .vdd(vdd), .A(_11163_), .Y(_11167_) );
AOI21X1 AOI21X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_11165_), .B(_11166_), .C(_11167_), .Y(_11168_) );
OAI21X1 OAI21X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_11164_), .B(_11168_), .C(_11088_), .Y(_11170_) );
NAND3X1 NAND3X1_2509 ( .gnd(gnd), .vdd(vdd), .A(_11167_), .B(_11165_), .C(_11166_), .Y(_11171_) );
OAI21X1 OAI21X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_11157_), .B(_11162_), .C(_11163_), .Y(_11172_) );
NAND3X1 NAND3X1_2510 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf1_), .B(_11171_), .C(_11172_), .Y(_11173_) );
NAND3X1 NAND3X1_2511 ( .gnd(gnd), .vdd(vdd), .A(_11087_), .B(_11173_), .C(_11170_), .Y(_11174_) );
AOI21X1 AOI21X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_11171_), .B(_11172_), .C(bloque_datos_45_bF_buf0_), .Y(_11175_) );
NOR3X1 NOR3X1_325 ( .gnd(gnd), .vdd(vdd), .A(_11168_), .B(_11088_), .C(_11164_), .Y(_11176_) );
OAI21X1 OAI21X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_11176_), .B(_11175_), .C(_10795_), .Y(_11177_) );
NAND3X1 NAND3X1_2512 ( .gnd(gnd), .vdd(vdd), .A(_11174_), .B(_11177_), .C(_11086_), .Y(_11178_) );
OAI21X1 OAI21X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_10717_), .B(_10803_), .C(_10808_), .Y(_11179_) );
NAND3X1 NAND3X1_2513 ( .gnd(gnd), .vdd(vdd), .A(_10795_), .B(_11173_), .C(_11170_), .Y(_11181_) );
OAI21X1 OAI21X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_11176_), .B(_11175_), .C(_11087_), .Y(_11182_) );
NAND3X1 NAND3X1_2514 ( .gnd(gnd), .vdd(vdd), .A(_11181_), .B(_11179_), .C(_11182_), .Y(_11183_) );
XOR2X1 XOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_9127_), .B(_11641_), .Y(_11184_) );
INVX1 INVX1_1529 ( .gnd(gnd), .vdd(vdd), .A(_11184_), .Y(_11185_) );
NAND3X1 NAND3X1_2515 ( .gnd(gnd), .vdd(vdd), .A(_11185_), .B(_11183_), .C(_11178_), .Y(_11186_) );
AOI21X1 AOI21X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_11181_), .B(_11182_), .C(_11179_), .Y(_11187_) );
AOI21X1 AOI21X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_11174_), .B(_11177_), .C(_11086_), .Y(_11188_) );
OAI21X1 OAI21X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_11188_), .B(_11187_), .C(_11184_), .Y(_11189_) );
NAND3X1 NAND3X1_2516 ( .gnd(gnd), .vdd(vdd), .A(_11085_), .B(_11186_), .C(_11189_), .Y(_11190_) );
NAND3X1 NAND3X1_2517 ( .gnd(gnd), .vdd(vdd), .A(_11184_), .B(_11183_), .C(_11178_), .Y(_11192_) );
OAI21X1 OAI21X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_11188_), .B(_11187_), .C(_11185_), .Y(_11193_) );
NAND3X1 NAND3X1_2518 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf1_), .B(_11192_), .C(_11193_), .Y(_11194_) );
NAND3X1 NAND3X1_2519 ( .gnd(gnd), .vdd(vdd), .A(_11084_), .B(_11190_), .C(_11194_), .Y(_11195_) );
AOI21X1 AOI21X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_11192_), .B(_11193_), .C(bloque_datos_61_bF_buf0_), .Y(_11196_) );
AOI21X1 AOI21X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_11186_), .B(_11189_), .C(_11085_), .Y(_11197_) );
OAI21X1 OAI21X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_11196_), .B(_11197_), .C(_10824_), .Y(_11198_) );
NAND3X1 NAND3X1_2520 ( .gnd(gnd), .vdd(vdd), .A(_11195_), .B(_11198_), .C(_11083_), .Y(_11199_) );
OAI21X1 OAI21X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_10830_), .B(_10832_), .C(_10822_), .Y(_11200_) );
NAND3X1 NAND3X1_2521 ( .gnd(gnd), .vdd(vdd), .A(_10824_), .B(_11190_), .C(_11194_), .Y(_11201_) );
OAI21X1 OAI21X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_11196_), .B(_11197_), .C(_11084_), .Y(_11203_) );
NAND3X1 NAND3X1_2522 ( .gnd(gnd), .vdd(vdd), .A(_11201_), .B(_11200_), .C(_11203_), .Y(_11204_) );
XNOR2X1 XNOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_9132_), .B(_11707_), .Y(_11205_) );
INVX1 INVX1_1530 ( .gnd(gnd), .vdd(vdd), .A(_11205_), .Y(_11206_) );
NAND3X1 NAND3X1_2523 ( .gnd(gnd), .vdd(vdd), .A(_11206_), .B(_11204_), .C(_11199_), .Y(_11207_) );
AOI21X1 AOI21X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_11201_), .B(_11203_), .C(_11200_), .Y(_11208_) );
AOI21X1 AOI21X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_11195_), .B(_11198_), .C(_11083_), .Y(_11209_) );
OAI21X1 OAI21X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_11208_), .B(_11209_), .C(_11205_), .Y(_11210_) );
NAND3X1 NAND3X1_2524 ( .gnd(gnd), .vdd(vdd), .A(_11082_), .B(_11207_), .C(_11210_), .Y(_11211_) );
NAND3X1 NAND3X1_2525 ( .gnd(gnd), .vdd(vdd), .A(_11205_), .B(_11204_), .C(_11199_), .Y(_11212_) );
OAI21X1 OAI21X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_11208_), .B(_11209_), .C(_11206_), .Y(_11214_) );
NAND3X1 NAND3X1_2526 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf1_), .B(_11212_), .C(_11214_), .Y(_11215_) );
NAND3X1 NAND3X1_2527 ( .gnd(gnd), .vdd(vdd), .A(_11080_), .B(_11211_), .C(_11215_), .Y(_11216_) );
AOI21X1 AOI21X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_11212_), .B(_11214_), .C(bloque_datos_77_bF_buf0_), .Y(_11217_) );
AOI21X1 AOI21X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_11207_), .B(_11210_), .C(_11082_), .Y(_11218_) );
OAI21X1 OAI21X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_11217_), .B(_11218_), .C(_10847_), .Y(_11219_) );
NAND3X1 NAND3X1_2528 ( .gnd(gnd), .vdd(vdd), .A(_11216_), .B(_11219_), .C(_11079_), .Y(_11220_) );
OAI21X1 OAI21X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_10855_), .B(_10853_), .C(_10845_), .Y(_11221_) );
NAND3X1 NAND3X1_2529 ( .gnd(gnd), .vdd(vdd), .A(_10847_), .B(_11211_), .C(_11215_), .Y(_11222_) );
OAI21X1 OAI21X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_11217_), .B(_11218_), .C(_11080_), .Y(_11223_) );
NAND3X1 NAND3X1_2530 ( .gnd(gnd), .vdd(vdd), .A(_11222_), .B(_11221_), .C(_11223_), .Y(_11225_) );
XNOR2X1 XNOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_9138_), .B(_11751_), .Y(_11226_) );
INVX1 INVX1_1531 ( .gnd(gnd), .vdd(vdd), .A(_11226_), .Y(_11227_) );
NAND3X1 NAND3X1_2531 ( .gnd(gnd), .vdd(vdd), .A(_11227_), .B(_11225_), .C(_11220_), .Y(_11228_) );
AOI21X1 AOI21X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_11222_), .B(_11223_), .C(_11221_), .Y(_11229_) );
AOI21X1 AOI21X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_11216_), .B(_11219_), .C(_11079_), .Y(_11230_) );
OAI21X1 OAI21X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_11229_), .B(_11230_), .C(_11226_), .Y(_11231_) );
NAND3X1 NAND3X1_2532 ( .gnd(gnd), .vdd(vdd), .A(_11078_), .B(_11228_), .C(_11231_), .Y(_11232_) );
NOR3X1 NOR3X1_326 ( .gnd(gnd), .vdd(vdd), .A(_11229_), .B(_11226_), .C(_11230_), .Y(_11233_) );
AOI21X1 AOI21X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_11225_), .B(_11220_), .C(_11227_), .Y(_11234_) );
OAI21X1 OAI21X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_11233_), .B(_11234_), .C(bloque_datos_93_bF_buf2_), .Y(_11236_) );
NAND3X1 NAND3X1_2533 ( .gnd(gnd), .vdd(vdd), .A(_10863_), .B(_11232_), .C(_11236_), .Y(_11237_) );
INVX1 INVX1_1532 ( .gnd(gnd), .vdd(vdd), .A(_10863_), .Y(_11238_) );
NOR3X1 NOR3X1_327 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf1_), .B(_11234_), .C(_11233_), .Y(_11239_) );
AOI21X1 AOI21X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_11228_), .B(_11231_), .C(_11078_), .Y(_11240_) );
OAI21X1 OAI21X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_11239_), .B(_11240_), .C(_11238_), .Y(_11241_) );
AOI21X1 AOI21X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_11237_), .B(_11241_), .C(_11077_), .Y(_11242_) );
AOI21X1 AOI21X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_10872_), .B(_10875_), .C(_10867_), .Y(_11243_) );
NAND3X1 NAND3X1_2534 ( .gnd(gnd), .vdd(vdd), .A(_11238_), .B(_11232_), .C(_11236_), .Y(_11244_) );
OAI21X1 OAI21X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_11239_), .B(_11240_), .C(_10863_), .Y(_11245_) );
AOI21X1 AOI21X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_11244_), .B(_11245_), .C(_11243_), .Y(_11247_) );
OAI21X1 OAI21X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_11242_), .B(_11247_), .C(_11849_), .Y(_11248_) );
NAND3X1 NAND3X1_2535 ( .gnd(gnd), .vdd(vdd), .A(_11243_), .B(_11244_), .C(_11245_), .Y(_11249_) );
NAND3X1 NAND3X1_2536 ( .gnd(gnd), .vdd(vdd), .A(_11077_), .B(_11237_), .C(_11241_), .Y(_11250_) );
NAND3X1 NAND3X1_2537 ( .gnd(gnd), .vdd(vdd), .A(_11860_), .B(_11249_), .C(_11250_), .Y(_11251_) );
NAND2X1 NAND2X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_11251_), .B(_11248_), .Y(_11252_) );
NAND3X1 NAND3X1_2538 ( .gnd(gnd), .vdd(vdd), .A(_11076_), .B(_9145_), .C(_11252_), .Y(_11253_) );
OAI21X1 OAI21X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_11242_), .B(_11247_), .C(_11860_), .Y(_11254_) );
NAND3X1 NAND3X1_2539 ( .gnd(gnd), .vdd(vdd), .A(_11849_), .B(_11249_), .C(_11250_), .Y(_11255_) );
NAND3X1 NAND3X1_2540 ( .gnd(gnd), .vdd(vdd), .A(_9145_), .B(_11255_), .C(_11254_), .Y(_11256_) );
NAND2X1 NAND2X1_1442 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_141_), .B(_11256_), .Y(_11258_) );
AOI21X1 AOI21X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_11253_), .B(_11258_), .C(_10891_), .Y(_11259_) );
INVX1 INVX1_1533 ( .gnd(gnd), .vdd(vdd), .A(_10891_), .Y(_11260_) );
NAND3X1 NAND3X1_2541 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_141_), .B(_9145_), .C(_11252_), .Y(_11261_) );
NAND2X1 NAND2X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_11076_), .B(_11256_), .Y(_11262_) );
AOI21X1 AOI21X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_11261_), .B(_11262_), .C(_11260_), .Y(_11263_) );
OAI21X1 OAI21X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_11259_), .B(_11263_), .C(_11075_), .Y(_11264_) );
OAI21X1 OAI21X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_10703_), .B(_10893_), .C(_10896_), .Y(_11265_) );
NAND3X1 NAND3X1_2542 ( .gnd(gnd), .vdd(vdd), .A(_11260_), .B(_11261_), .C(_11262_), .Y(_11266_) );
NAND3X1 NAND3X1_2543 ( .gnd(gnd), .vdd(vdd), .A(_10891_), .B(_11253_), .C(_11258_), .Y(_11267_) );
NAND3X1 NAND3X1_2544 ( .gnd(gnd), .vdd(vdd), .A(_11266_), .B(_11267_), .C(_11265_), .Y(_11269_) );
NAND3X1 NAND3X1_2545 ( .gnd(gnd), .vdd(vdd), .A(_11074_), .B(_11269_), .C(_11264_), .Y(_11270_) );
AOI21X1 AOI21X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_11266_), .B(_11267_), .C(_11265_), .Y(_11271_) );
NOR3X1 NOR3X1_328 ( .gnd(gnd), .vdd(vdd), .A(_11259_), .B(_11075_), .C(_11263_), .Y(_11272_) );
OAI21X1 OAI21X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_11272_), .B(_11271_), .C(_11926_), .Y(_11273_) );
NAND2X1 NAND2X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_11270_), .B(_11273_), .Y(_11274_) );
NAND3X1 NAND3X1_2546 ( .gnd(gnd), .vdd(vdd), .A(_11073_), .B(_9153_), .C(_11274_), .Y(_11275_) );
OAI21X1 OAI21X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_11272_), .B(_11271_), .C(_11074_), .Y(_11276_) );
NAND3X1 NAND3X1_2547 ( .gnd(gnd), .vdd(vdd), .A(_11926_), .B(_11269_), .C(_11264_), .Y(_11277_) );
NAND3X1 NAND3X1_2548 ( .gnd(gnd), .vdd(vdd), .A(_9153_), .B(_11277_), .C(_11276_), .Y(_11278_) );
NAND2X1 NAND2X1_1445 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_157_), .B(_11278_), .Y(_11280_) );
AOI21X1 AOI21X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_11275_), .B(_11280_), .C(_10911_), .Y(_11281_) );
INVX1 INVX1_1534 ( .gnd(gnd), .vdd(vdd), .A(_10911_), .Y(_11282_) );
NAND3X1 NAND3X1_2549 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_157_), .B(_9153_), .C(_11274_), .Y(_11283_) );
NAND2X1 NAND2X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_11073_), .B(_11278_), .Y(_11284_) );
AOI21X1 AOI21X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_11283_), .B(_11284_), .C(_11282_), .Y(_11285_) );
OAI21X1 OAI21X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_11281_), .B(_11285_), .C(_11072_), .Y(_11286_) );
OAI21X1 OAI21X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_10913_), .B(_10701_), .C(_10918_), .Y(_11287_) );
NAND3X1 NAND3X1_2550 ( .gnd(gnd), .vdd(vdd), .A(_11282_), .B(_11283_), .C(_11284_), .Y(_11288_) );
NAND3X1 NAND3X1_2551 ( .gnd(gnd), .vdd(vdd), .A(_10911_), .B(_11275_), .C(_11280_), .Y(_11289_) );
NAND3X1 NAND3X1_2552 ( .gnd(gnd), .vdd(vdd), .A(_11288_), .B(_11289_), .C(_11287_), .Y(_11291_) );
NAND3X1 NAND3X1_2553 ( .gnd(gnd), .vdd(vdd), .A(_11071_), .B(_11291_), .C(_11286_), .Y(_11292_) );
AOI21X1 AOI21X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_11288_), .B(_11289_), .C(_11287_), .Y(_11293_) );
NOR3X1 NOR3X1_329 ( .gnd(gnd), .vdd(vdd), .A(_11281_), .B(_11072_), .C(_11285_), .Y(_11294_) );
OAI21X1 OAI21X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_11294_), .B(_11293_), .C(_12010_), .Y(_11295_) );
NAND2X1 NAND2X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_11292_), .B(_11295_), .Y(_11296_) );
NAND3X1 NAND3X1_2554 ( .gnd(gnd), .vdd(vdd), .A(_11069_), .B(_9161_), .C(_11296_), .Y(_11297_) );
OAI21X1 OAI21X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_11294_), .B(_11293_), .C(_11071_), .Y(_11298_) );
NAND3X1 NAND3X1_2555 ( .gnd(gnd), .vdd(vdd), .A(_12010_), .B(_11291_), .C(_11286_), .Y(_11299_) );
NAND3X1 NAND3X1_2556 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .B(_11299_), .C(_11298_), .Y(_11300_) );
NAND2X1 NAND2X1_1448 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_173_), .B(_11300_), .Y(_11302_) );
AOI21X1 AOI21X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_11297_), .B(_11302_), .C(_10924_), .Y(_11303_) );
INVX1 INVX1_1535 ( .gnd(gnd), .vdd(vdd), .A(_10924_), .Y(_11304_) );
NAND3X1 NAND3X1_2557 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_173_), .B(_9161_), .C(_11296_), .Y(_11305_) );
NAND2X1 NAND2X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_11069_), .B(_11300_), .Y(_11306_) );
AOI21X1 AOI21X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_11305_), .B(_11306_), .C(_11304_), .Y(_11307_) );
OAI21X1 OAI21X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_11303_), .B(_11307_), .C(_11068_), .Y(_11308_) );
OAI21X1 OAI21X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_10940_), .B(_10942_), .C(_10933_), .Y(_11309_) );
NAND3X1 NAND3X1_2558 ( .gnd(gnd), .vdd(vdd), .A(_11304_), .B(_11305_), .C(_11306_), .Y(_11310_) );
NAND3X1 NAND3X1_2559 ( .gnd(gnd), .vdd(vdd), .A(_10924_), .B(_11297_), .C(_11302_), .Y(_11311_) );
NAND3X1 NAND3X1_2560 ( .gnd(gnd), .vdd(vdd), .A(_11310_), .B(_11311_), .C(_11309_), .Y(_11313_) );
NAND3X1 NAND3X1_2561 ( .gnd(gnd), .vdd(vdd), .A(_12019_), .B(_11313_), .C(_11308_), .Y(_11314_) );
AOI21X1 AOI21X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_11310_), .B(_11311_), .C(_11309_), .Y(_11315_) );
NOR3X1 NOR3X1_330 ( .gnd(gnd), .vdd(vdd), .A(_11303_), .B(_11068_), .C(_11307_), .Y(_11316_) );
OAI21X1 OAI21X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_11316_), .B(_11315_), .C(_12018_), .Y(_11317_) );
NAND2X1 NAND2X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_11314_), .B(_11317_), .Y(_11318_) );
NAND3X1 NAND3X1_2562 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_189_), .B(_9169_), .C(_11318_), .Y(_11319_) );
INVX1 INVX1_1536 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_189_), .Y(_11320_) );
OAI21X1 OAI21X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_11316_), .B(_11315_), .C(_12019_), .Y(_11321_) );
NAND3X1 NAND3X1_2563 ( .gnd(gnd), .vdd(vdd), .A(_12018_), .B(_11313_), .C(_11308_), .Y(_11322_) );
NAND3X1 NAND3X1_2564 ( .gnd(gnd), .vdd(vdd), .A(_9169_), .B(_11322_), .C(_11321_), .Y(_11324_) );
NAND2X1 NAND2X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_11320_), .B(_11324_), .Y(_11325_) );
NAND3X1 NAND3X1_2565 ( .gnd(gnd), .vdd(vdd), .A(_11067_), .B(_11319_), .C(_11325_), .Y(_11326_) );
NAND3X1 NAND3X1_2566 ( .gnd(gnd), .vdd(vdd), .A(_11320_), .B(_9169_), .C(_11318_), .Y(_11327_) );
NAND2X1 NAND2X1_1452 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_189_), .B(_11324_), .Y(_11328_) );
NAND3X1 NAND3X1_2567 ( .gnd(gnd), .vdd(vdd), .A(_10949_), .B(_11327_), .C(_11328_), .Y(_11329_) );
AOI21X1 AOI21X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_11326_), .B(_11329_), .C(_11066_), .Y(_11330_) );
AOI21X1 AOI21X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_10694_), .B(_10959_), .C(_10964_), .Y(_11331_) );
AOI21X1 AOI21X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_11327_), .B(_11328_), .C(_10949_), .Y(_11332_) );
AOI21X1 AOI21X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_11319_), .B(_11325_), .C(_11067_), .Y(_11333_) );
NOR3X1 NOR3X1_331 ( .gnd(gnd), .vdd(vdd), .A(_11332_), .B(_11331_), .C(_11333_), .Y(_11335_) );
OAI21X1 OAI21X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_11335_), .B(_11330_), .C(_12027_), .Y(_11336_) );
INVX1 INVX1_1537 ( .gnd(gnd), .vdd(vdd), .A(_12027_), .Y(_11337_) );
OAI21X1 OAI21X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_11332_), .B(_11333_), .C(_11331_), .Y(_11338_) );
NAND3X1 NAND3X1_2568 ( .gnd(gnd), .vdd(vdd), .A(_11326_), .B(_11329_), .C(_11066_), .Y(_11339_) );
NAND3X1 NAND3X1_2569 ( .gnd(gnd), .vdd(vdd), .A(_11337_), .B(_11338_), .C(_11339_), .Y(_11340_) );
NAND2X1 NAND2X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_11340_), .B(_11336_), .Y(_11341_) );
NAND3X1 NAND3X1_2570 ( .gnd(gnd), .vdd(vdd), .A(_11065_), .B(_9177_), .C(_11341_), .Y(_11342_) );
OAI21X1 OAI21X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_11335_), .B(_11330_), .C(_11337_), .Y(_11343_) );
NAND3X1 NAND3X1_2571 ( .gnd(gnd), .vdd(vdd), .A(_12027_), .B(_11338_), .C(_11339_), .Y(_11344_) );
NAND3X1 NAND3X1_2572 ( .gnd(gnd), .vdd(vdd), .A(_9177_), .B(_11344_), .C(_11343_), .Y(_11346_) );
NAND2X1 NAND2X1_1454 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_205_), .B(_11346_), .Y(_11347_) );
AOI21X1 AOI21X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_11342_), .B(_11347_), .C(_10980_), .Y(_11348_) );
INVX1 INVX1_1538 ( .gnd(gnd), .vdd(vdd), .A(_10980_), .Y(_11349_) );
NAND3X1 NAND3X1_2573 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_205_), .B(_9177_), .C(_11341_), .Y(_11350_) );
NAND2X1 NAND2X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_11065_), .B(_11346_), .Y(_11351_) );
AOI21X1 AOI21X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_11350_), .B(_11351_), .C(_11349_), .Y(_11352_) );
OAI21X1 OAI21X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_11348_), .B(_11352_), .C(_11064_), .Y(_11353_) );
OAI21X1 OAI21X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_10982_), .B(_10693_), .C(_10987_), .Y(_11354_) );
NAND3X1 NAND3X1_2574 ( .gnd(gnd), .vdd(vdd), .A(_11349_), .B(_11350_), .C(_11351_), .Y(_11355_) );
NAND3X1 NAND3X1_2575 ( .gnd(gnd), .vdd(vdd), .A(_10980_), .B(_11342_), .C(_11347_), .Y(_11357_) );
NAND3X1 NAND3X1_2576 ( .gnd(gnd), .vdd(vdd), .A(_11355_), .B(_11357_), .C(_11354_), .Y(_11358_) );
NAND3X1 NAND3X1_2577 ( .gnd(gnd), .vdd(vdd), .A(_12035_), .B(_11358_), .C(_11353_), .Y(_11359_) );
NAND2X1 NAND2X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_11358_), .B(_11353_), .Y(_11360_) );
AOI21X1 AOI21X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_12036_), .B(_11360_), .C(_9186_), .Y(_11361_) );
NAND3X1 NAND3X1_2578 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_221_), .B(_11359_), .C(_11361_), .Y(_11362_) );
INVX1 INVX1_1539 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_221_), .Y(_11363_) );
AOI21X1 AOI21X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_11355_), .B(_11357_), .C(_11354_), .Y(_11364_) );
NOR3X1 NOR3X1_332 ( .gnd(gnd), .vdd(vdd), .A(_11064_), .B(_11348_), .C(_11352_), .Y(_11365_) );
OAI21X1 OAI21X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_11365_), .B(_11364_), .C(_12036_), .Y(_11366_) );
NAND3X1 NAND3X1_2579 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_11359_), .C(_11366_), .Y(_11368_) );
NAND2X1 NAND2X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_11363_), .B(_11368_), .Y(_11369_) );
NAND3X1 NAND3X1_2580 ( .gnd(gnd), .vdd(vdd), .A(_11063_), .B(_11362_), .C(_11369_), .Y(_11370_) );
NAND3X1 NAND3X1_2581 ( .gnd(gnd), .vdd(vdd), .A(_11363_), .B(_11359_), .C(_11361_), .Y(_11371_) );
NAND2X1 NAND2X1_1458 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_221_), .B(_11368_), .Y(_11372_) );
NAND3X1 NAND3X1_2582 ( .gnd(gnd), .vdd(vdd), .A(_11003_), .B(_11371_), .C(_11372_), .Y(_11373_) );
AOI21X1 AOI21X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_11370_), .B(_11373_), .C(_11062_), .Y(_11374_) );
AOI21X1 AOI21X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_11010_), .B(_11012_), .C(_11002_), .Y(_11375_) );
AOI21X1 AOI21X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_11371_), .B(_11372_), .C(_11003_), .Y(_11376_) );
AOI21X1 AOI21X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_11362_), .B(_11369_), .C(_11063_), .Y(_11377_) );
NOR3X1 NOR3X1_333 ( .gnd(gnd), .vdd(vdd), .A(_11376_), .B(_11375_), .C(_11377_), .Y(_11379_) );
OAI21X1 OAI21X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_11379_), .B(_11374_), .C(_12044_), .Y(_11380_) );
INVX1 INVX1_1540 ( .gnd(gnd), .vdd(vdd), .A(_12044_), .Y(_11381_) );
OAI21X1 OAI21X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_11376_), .B(_11377_), .C(_11375_), .Y(_11382_) );
NAND3X1 NAND3X1_2583 ( .gnd(gnd), .vdd(vdd), .A(_11370_), .B(_11373_), .C(_11062_), .Y(_11383_) );
NAND3X1 NAND3X1_2584 ( .gnd(gnd), .vdd(vdd), .A(_11381_), .B(_11383_), .C(_11382_), .Y(_11384_) );
NAND2X1 NAND2X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_11384_), .B(_11380_), .Y(_11385_) );
NAND3X1 NAND3X1_2585 ( .gnd(gnd), .vdd(vdd), .A(_11061_), .B(_9193_), .C(_11385_), .Y(_11386_) );
OAI21X1 OAI21X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_11379_), .B(_11374_), .C(_11381_), .Y(_11387_) );
NAND3X1 NAND3X1_2586 ( .gnd(gnd), .vdd(vdd), .A(_12044_), .B(_11383_), .C(_11382_), .Y(_11388_) );
NAND3X1 NAND3X1_2587 ( .gnd(gnd), .vdd(vdd), .A(_9193_), .B(_11388_), .C(_11387_), .Y(_11390_) );
NAND2X1 NAND2X1_1460 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_237_), .B(_11390_), .Y(_11391_) );
AOI21X1 AOI21X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_11386_), .B(_11391_), .C(_11018_), .Y(_11392_) );
INVX1 INVX1_1541 ( .gnd(gnd), .vdd(vdd), .A(_11018_), .Y(_11393_) );
NAND3X1 NAND3X1_2588 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_237_), .B(_9193_), .C(_11385_), .Y(_11394_) );
NAND2X1 NAND2X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_11061_), .B(_11390_), .Y(_11395_) );
AOI21X1 AOI21X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_11394_), .B(_11395_), .C(_11393_), .Y(_11396_) );
OAI21X1 OAI21X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_11392_), .B(_11396_), .C(_11060_), .Y(_11397_) );
OAI21X1 OAI21X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_11033_), .B(_11040_), .C(_11026_), .Y(_11398_) );
NAND3X1 NAND3X1_2589 ( .gnd(gnd), .vdd(vdd), .A(_11393_), .B(_11394_), .C(_11395_), .Y(_11399_) );
NAND3X1 NAND3X1_2590 ( .gnd(gnd), .vdd(vdd), .A(_11018_), .B(_11386_), .C(_11391_), .Y(_11401_) );
NAND3X1 NAND3X1_2591 ( .gnd(gnd), .vdd(vdd), .A(_11399_), .B(_11401_), .C(_11398_), .Y(_11402_) );
NAND3X1 NAND3X1_2592 ( .gnd(gnd), .vdd(vdd), .A(_12241_), .B(_11397_), .C(_11402_), .Y(_11403_) );
AOI21X1 AOI21X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_11399_), .B(_11401_), .C(_11398_), .Y(_11404_) );
NOR3X1 NOR3X1_334 ( .gnd(gnd), .vdd(vdd), .A(_11392_), .B(_11060_), .C(_11396_), .Y(_11405_) );
OAI21X1 OAI21X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_11405_), .B(_11404_), .C(_12052_), .Y(_11406_) );
NAND2X1 NAND2X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_11403_), .B(_11406_), .Y(_11407_) );
NAND3X1 NAND3X1_2593 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_253_), .B(_9201_), .C(_11407_), .Y(_11408_) );
INVX1 INVX1_1542 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_253_), .Y(_11409_) );
OAI21X1 OAI21X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_11405_), .B(_11404_), .C(_12241_), .Y(_11410_) );
NAND3X1 NAND3X1_2594 ( .gnd(gnd), .vdd(vdd), .A(_12052_), .B(_11397_), .C(_11402_), .Y(_11412_) );
NAND3X1 NAND3X1_2595 ( .gnd(gnd), .vdd(vdd), .A(_9201_), .B(_11412_), .C(_11410_), .Y(_11413_) );
NAND2X1 NAND2X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_11409_), .B(_11413_), .Y(_11414_) );
NAND3X1 NAND3X1_2596 ( .gnd(gnd), .vdd(vdd), .A(_11058_), .B(_11408_), .C(_11414_), .Y(_11415_) );
INVX1 INVX1_1543 ( .gnd(gnd), .vdd(vdd), .A(_11058_), .Y(_11416_) );
NAND2X1 NAND2X1_1464 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_253_), .B(_11413_), .Y(_11417_) );
OR2X2 OR2X2_254 ( .gnd(gnd), .vdd(vdd), .A(_11413_), .B(module_2_W_253_), .Y(_11418_) );
NAND3X1 NAND3X1_2597 ( .gnd(gnd), .vdd(vdd), .A(_11416_), .B(_11417_), .C(_11418_), .Y(_11419_) );
NAND2X1 NAND2X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_11415_), .B(_11419_), .Y(_11420_) );
XNOR2X1 XNOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_11420_), .B(_11056_), .Y(module_2_H_21_) );
AOI21X1 AOI21X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_11408_), .B(_11414_), .C(_11058_), .Y(_11422_) );
AOI21X1 AOI21X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_11056_), .B(_11415_), .C(_11422_), .Y(_11423_) );
INVX1 INVX1_1544 ( .gnd(gnd), .vdd(vdd), .A(_11423_), .Y(_11424_) );
INVX1 INVX1_1545 ( .gnd(gnd), .vdd(vdd), .A(_11417_), .Y(_11425_) );
OAI21X1 OAI21X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_11396_), .B(_11060_), .C(_11399_), .Y(_11426_) );
OAI21X1 OAI21X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_11377_), .B(_11375_), .C(_11370_), .Y(_11427_) );
OAI21X1 OAI21X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_11064_), .B(_11352_), .C(_11355_), .Y(_11428_) );
OAI21X1 OAI21X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_11333_), .B(_11331_), .C(_11326_), .Y(_11429_) );
INVX1 INVX1_1546 ( .gnd(gnd), .vdd(vdd), .A(_11429_), .Y(_11430_) );
INVX1 INVX1_1547 ( .gnd(gnd), .vdd(vdd), .A(_11327_), .Y(_11431_) );
OAI21X1 OAI21X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_11307_), .B(_11068_), .C(_11310_), .Y(_11433_) );
INVX1 INVX1_1548 ( .gnd(gnd), .vdd(vdd), .A(_11433_), .Y(_11434_) );
INVX1 INVX1_1549 ( .gnd(gnd), .vdd(vdd), .A(_11297_), .Y(_11435_) );
OAI21X1 OAI21X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_11285_), .B(_11072_), .C(_11288_), .Y(_11436_) );
INVX1 INVX1_1550 ( .gnd(gnd), .vdd(vdd), .A(_11436_), .Y(_11437_) );
INVX1 INVX1_1551 ( .gnd(gnd), .vdd(vdd), .A(_11275_), .Y(_11438_) );
OAI21X1 OAI21X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_11263_), .B(_11075_), .C(_11266_), .Y(_11439_) );
NAND2X1 NAND2X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_11237_), .B(_11250_), .Y(_11440_) );
INVX1 INVX1_1552 ( .gnd(gnd), .vdd(vdd), .A(_11440_), .Y(_11441_) );
NAND2X1 NAND2X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_11222_), .B(_11225_), .Y(_11442_) );
NAND2X1 NAND2X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_11201_), .B(_11204_), .Y(_11444_) );
NAND2X1 NAND2X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_11181_), .B(_11183_), .Y(_11445_) );
NAND2X1 NAND2X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_11152_), .B(_11166_), .Y(_11446_) );
NAND2X1 NAND2X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_11138_), .B(_11140_), .Y(_11447_) );
OAI21X1 OAI21X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_11116_), .B(_11117_), .C(_11113_), .Y(_11448_) );
INVX1 INVX1_1553 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_30_), .Y(_11449_) );
NOR2X1 NOR2X1_852 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_12_), .B(module_2_W_13_), .Y(_11450_) );
XNOR2X1 XNOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_11450_), .B(module_2_W_14_), .Y(_11451_) );
XNOR2X1 XNOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_9591_), .B(module_2_W_10_), .Y(_11452_) );
XNOR2X1 XNOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_11452_), .B(_11451_), .Y(_11453_) );
OR2X2 OR2X2_255 ( .gnd(gnd), .vdd(vdd), .A(_11453_), .B(_11449_), .Y(_11455_) );
NAND2X1 NAND2X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_11449_), .B(_11453_), .Y(_11456_) );
NAND2X1 NAND2X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_11456_), .B(_11455_), .Y(_11457_) );
XNOR2X1 XNOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_11457_), .B(_11109_), .Y(_11458_) );
XOR2X1 XOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_11458_), .B(_11448_), .Y(_11459_) );
XNOR2X1 XNOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_9615_), .B(_9650_), .Y(_11460_) );
XOR2X1 XOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_11459_), .B(_11460_), .Y(_11461_) );
NAND2X1 NAND2X1_1474 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf3_), .B(_11461_), .Y(_11462_) );
INVX1 INVX1_1554 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf2_), .Y(_11463_) );
XNOR2X1 XNOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_11459_), .B(_11460_), .Y(_11464_) );
NAND2X1 NAND2X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_11463_), .B(_11464_), .Y(_11466_) );
NAND3X1 NAND3X1_2598 ( .gnd(gnd), .vdd(vdd), .A(_11133_), .B(_11466_), .C(_11462_), .Y(_11467_) );
NAND2X1 NAND2X1_1476 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf1_), .B(_11464_), .Y(_11468_) );
NAND2X1 NAND2X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_11463_), .B(_11461_), .Y(_11469_) );
NAND3X1 NAND3X1_2599 ( .gnd(gnd), .vdd(vdd), .A(_11130_), .B(_11468_), .C(_11469_), .Y(_11470_) );
NAND3X1 NAND3X1_2600 ( .gnd(gnd), .vdd(vdd), .A(_11447_), .B(_11467_), .C(_11470_), .Y(_11471_) );
AOI21X1 AOI21X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_11467_), .B(_11470_), .C(_11447_), .Y(_11472_) );
INVX1 INVX1_1555 ( .gnd(gnd), .vdd(vdd), .A(_11472_), .Y(_11473_) );
XNOR2X1 XNOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_9685_), .B(_9636_), .Y(_11474_) );
NAND3X1 NAND3X1_2601 ( .gnd(gnd), .vdd(vdd), .A(_11471_), .B(_11474_), .C(_11473_), .Y(_11475_) );
INVX1 INVX1_1556 ( .gnd(gnd), .vdd(vdd), .A(_11471_), .Y(_11477_) );
INVX1 INVX1_1557 ( .gnd(gnd), .vdd(vdd), .A(_11474_), .Y(_11478_) );
OAI21X1 OAI21X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_11477_), .B(_11472_), .C(_11478_), .Y(_11479_) );
NAND3X1 NAND3X1_2602 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf1_), .B(_11475_), .C(_11479_), .Y(_11480_) );
INVX1 INVX1_1558 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf0_), .Y(_11481_) );
OAI21X1 OAI21X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_11477_), .B(_11472_), .C(_11474_), .Y(_11482_) );
NAND3X1 NAND3X1_2603 ( .gnd(gnd), .vdd(vdd), .A(_11471_), .B(_11478_), .C(_11473_), .Y(_11483_) );
NAND3X1 NAND3X1_2604 ( .gnd(gnd), .vdd(vdd), .A(_11481_), .B(_11483_), .C(_11482_), .Y(_11484_) );
NAND3X1 NAND3X1_2605 ( .gnd(gnd), .vdd(vdd), .A(_11155_), .B(_11480_), .C(_11484_), .Y(_11485_) );
NAND3X1 NAND3X1_2606 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf3_), .B(_11483_), .C(_11482_), .Y(_11486_) );
NAND3X1 NAND3X1_2607 ( .gnd(gnd), .vdd(vdd), .A(_11481_), .B(_11475_), .C(_11479_), .Y(_11488_) );
NAND3X1 NAND3X1_2608 ( .gnd(gnd), .vdd(vdd), .A(_11151_), .B(_11486_), .C(_11488_), .Y(_11489_) );
NAND3X1 NAND3X1_2609 ( .gnd(gnd), .vdd(vdd), .A(_11446_), .B(_11485_), .C(_11489_), .Y(_11490_) );
INVX1 INVX1_1559 ( .gnd(gnd), .vdd(vdd), .A(_11446_), .Y(_11491_) );
NAND3X1 NAND3X1_2610 ( .gnd(gnd), .vdd(vdd), .A(_11155_), .B(_11486_), .C(_11488_), .Y(_11492_) );
NAND3X1 NAND3X1_2611 ( .gnd(gnd), .vdd(vdd), .A(_11151_), .B(_11480_), .C(_11484_), .Y(_11493_) );
NAND3X1 NAND3X1_2612 ( .gnd(gnd), .vdd(vdd), .A(_11491_), .B(_11492_), .C(_11493_), .Y(_11494_) );
XNOR2X1 XNOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_9723_), .B(_9673_), .Y(_11495_) );
NAND3X1 NAND3X1_2613 ( .gnd(gnd), .vdd(vdd), .A(_11495_), .B(_11490_), .C(_11494_), .Y(_11496_) );
AOI21X1 AOI21X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_11492_), .B(_11493_), .C(_11491_), .Y(_11497_) );
AOI21X1 AOI21X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_11485_), .B(_11489_), .C(_11446_), .Y(_11499_) );
INVX1 INVX1_1560 ( .gnd(gnd), .vdd(vdd), .A(_11495_), .Y(_11500_) );
OAI21X1 OAI21X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_11497_), .B(_11499_), .C(_11500_), .Y(_11501_) );
NAND3X1 NAND3X1_2614 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf2_), .B(_11496_), .C(_11501_), .Y(_11502_) );
INVX1 INVX1_1561 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf1_), .Y(_11503_) );
OAI21X1 OAI21X1_1830 ( .gnd(gnd), .vdd(vdd), .A(_11497_), .B(_11499_), .C(_11495_), .Y(_11504_) );
NAND3X1 NAND3X1_2615 ( .gnd(gnd), .vdd(vdd), .A(_11500_), .B(_11490_), .C(_11494_), .Y(_11505_) );
NAND3X1 NAND3X1_2616 ( .gnd(gnd), .vdd(vdd), .A(_11503_), .B(_11505_), .C(_11504_), .Y(_11506_) );
NAND3X1 NAND3X1_2617 ( .gnd(gnd), .vdd(vdd), .A(_11176_), .B(_11502_), .C(_11506_), .Y(_11507_) );
NAND3X1 NAND3X1_2618 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf0_), .B(_11505_), .C(_11504_), .Y(_11508_) );
NAND3X1 NAND3X1_2619 ( .gnd(gnd), .vdd(vdd), .A(_11503_), .B(_11496_), .C(_11501_), .Y(_11510_) );
NAND3X1 NAND3X1_2620 ( .gnd(gnd), .vdd(vdd), .A(_11173_), .B(_11508_), .C(_11510_), .Y(_11511_) );
NAND3X1 NAND3X1_2621 ( .gnd(gnd), .vdd(vdd), .A(_11445_), .B(_11507_), .C(_11511_), .Y(_11512_) );
INVX1 INVX1_1562 ( .gnd(gnd), .vdd(vdd), .A(_11445_), .Y(_11513_) );
NAND3X1 NAND3X1_2622 ( .gnd(gnd), .vdd(vdd), .A(_11176_), .B(_11508_), .C(_11510_), .Y(_11514_) );
NAND3X1 NAND3X1_2623 ( .gnd(gnd), .vdd(vdd), .A(_11173_), .B(_11502_), .C(_11506_), .Y(_11515_) );
NAND3X1 NAND3X1_2624 ( .gnd(gnd), .vdd(vdd), .A(_11513_), .B(_11514_), .C(_11515_), .Y(_11516_) );
XNOR2X1 XNOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_9762_), .B(_12339_), .Y(_11517_) );
NAND3X1 NAND3X1_2625 ( .gnd(gnd), .vdd(vdd), .A(_11517_), .B(_11512_), .C(_11516_), .Y(_11518_) );
AOI21X1 AOI21X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_11514_), .B(_11515_), .C(_11513_), .Y(_11519_) );
AOI21X1 AOI21X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_11507_), .B(_11511_), .C(_11445_), .Y(_11521_) );
INVX1 INVX1_1563 ( .gnd(gnd), .vdd(vdd), .A(_11517_), .Y(_11522_) );
OAI21X1 OAI21X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_11519_), .B(_11521_), .C(_11522_), .Y(_11523_) );
NAND3X1 NAND3X1_2626 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf1_), .B(_11518_), .C(_11523_), .Y(_11524_) );
INVX1 INVX1_1564 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf0_), .Y(_11525_) );
OAI21X1 OAI21X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_11519_), .B(_11521_), .C(_11517_), .Y(_11526_) );
NAND3X1 NAND3X1_2627 ( .gnd(gnd), .vdd(vdd), .A(_11522_), .B(_11512_), .C(_11516_), .Y(_11527_) );
NAND3X1 NAND3X1_2628 ( .gnd(gnd), .vdd(vdd), .A(_11525_), .B(_11527_), .C(_11526_), .Y(_11528_) );
NAND3X1 NAND3X1_2629 ( .gnd(gnd), .vdd(vdd), .A(_11197_), .B(_11524_), .C(_11528_), .Y(_11529_) );
NAND3X1 NAND3X1_2630 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf3_), .B(_11527_), .C(_11526_), .Y(_11530_) );
NAND3X1 NAND3X1_2631 ( .gnd(gnd), .vdd(vdd), .A(_11525_), .B(_11518_), .C(_11523_), .Y(_11532_) );
NAND3X1 NAND3X1_2632 ( .gnd(gnd), .vdd(vdd), .A(_11194_), .B(_11530_), .C(_11532_), .Y(_11533_) );
NAND3X1 NAND3X1_2633 ( .gnd(gnd), .vdd(vdd), .A(_11444_), .B(_11529_), .C(_11533_), .Y(_11534_) );
INVX2 INVX2_380 ( .gnd(gnd), .vdd(vdd), .A(_11444_), .Y(_11535_) );
AOI21X1 AOI21X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_11530_), .B(_11532_), .C(_11194_), .Y(_11536_) );
AOI21X1 AOI21X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_11524_), .B(_11528_), .C(_11197_), .Y(_11537_) );
OAI21X1 OAI21X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_11536_), .B(_11537_), .C(_11535_), .Y(_11538_) );
XOR2X1 XOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_9803_), .B(_9764_), .Y(_11539_) );
NAND3X1 NAND3X1_2634 ( .gnd(gnd), .vdd(vdd), .A(_11534_), .B(_11539_), .C(_11538_), .Y(_11540_) );
NOR3X1 NOR3X1_335 ( .gnd(gnd), .vdd(vdd), .A(_11536_), .B(_11535_), .C(_11537_), .Y(_11541_) );
AOI21X1 AOI21X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_11529_), .B(_11533_), .C(_11444_), .Y(_11543_) );
INVX1 INVX1_1565 ( .gnd(gnd), .vdd(vdd), .A(_11539_), .Y(_11544_) );
OAI21X1 OAI21X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_11541_), .B(_11543_), .C(_11544_), .Y(_11545_) );
NAND3X1 NAND3X1_2635 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf2_), .B(_11540_), .C(_11545_), .Y(_11546_) );
INVX1 INVX1_1566 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf1_), .Y(_11547_) );
OAI21X1 OAI21X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_11541_), .B(_11543_), .C(_11539_), .Y(_11548_) );
NAND3X1 NAND3X1_2636 ( .gnd(gnd), .vdd(vdd), .A(_11534_), .B(_11544_), .C(_11538_), .Y(_11549_) );
NAND3X1 NAND3X1_2637 ( .gnd(gnd), .vdd(vdd), .A(_11547_), .B(_11549_), .C(_11548_), .Y(_11550_) );
NAND3X1 NAND3X1_2638 ( .gnd(gnd), .vdd(vdd), .A(_11218_), .B(_11546_), .C(_11550_), .Y(_11551_) );
NAND3X1 NAND3X1_2639 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf0_), .B(_11549_), .C(_11548_), .Y(_11552_) );
NAND3X1 NAND3X1_2640 ( .gnd(gnd), .vdd(vdd), .A(_11547_), .B(_11540_), .C(_11545_), .Y(_11554_) );
NAND3X1 NAND3X1_2641 ( .gnd(gnd), .vdd(vdd), .A(_11215_), .B(_11552_), .C(_11554_), .Y(_11555_) );
NAND3X1 NAND3X1_2642 ( .gnd(gnd), .vdd(vdd), .A(_11442_), .B(_11551_), .C(_11555_), .Y(_11556_) );
INVX1 INVX1_1567 ( .gnd(gnd), .vdd(vdd), .A(_11442_), .Y(_11557_) );
NAND3X1 NAND3X1_2643 ( .gnd(gnd), .vdd(vdd), .A(_11218_), .B(_11552_), .C(_11554_), .Y(_11558_) );
NAND3X1 NAND3X1_2644 ( .gnd(gnd), .vdd(vdd), .A(_11215_), .B(_11546_), .C(_11550_), .Y(_11559_) );
NAND3X1 NAND3X1_2645 ( .gnd(gnd), .vdd(vdd), .A(_11557_), .B(_11558_), .C(_11559_), .Y(_11560_) );
XOR2X1 XOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_9843_), .B(_9805_), .Y(_11561_) );
INVX1 INVX1_1568 ( .gnd(gnd), .vdd(vdd), .A(_11561_), .Y(_11562_) );
NAND3X1 NAND3X1_2646 ( .gnd(gnd), .vdd(vdd), .A(_11562_), .B(_11556_), .C(_11560_), .Y(_11563_) );
AOI21X1 AOI21X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_11558_), .B(_11559_), .C(_11557_), .Y(_11565_) );
AOI21X1 AOI21X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_11551_), .B(_11555_), .C(_11442_), .Y(_11566_) );
OAI21X1 OAI21X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_11565_), .B(_11566_), .C(_11561_), .Y(_11567_) );
NAND3X1 NAND3X1_2647 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf3_), .B(_11563_), .C(_11567_), .Y(_11568_) );
INVX1 INVX1_1569 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf2_), .Y(_11569_) );
NAND3X1 NAND3X1_2648 ( .gnd(gnd), .vdd(vdd), .A(_11561_), .B(_11556_), .C(_11560_), .Y(_11570_) );
OAI21X1 OAI21X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_11565_), .B(_11566_), .C(_11562_), .Y(_11571_) );
NAND3X1 NAND3X1_2649 ( .gnd(gnd), .vdd(vdd), .A(_11569_), .B(_11570_), .C(_11571_), .Y(_11572_) );
NAND3X1 NAND3X1_2650 ( .gnd(gnd), .vdd(vdd), .A(_11240_), .B(_11568_), .C(_11572_), .Y(_11573_) );
NAND3X1 NAND3X1_2651 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf1_), .B(_11570_), .C(_11571_), .Y(_11574_) );
NAND3X1 NAND3X1_2652 ( .gnd(gnd), .vdd(vdd), .A(_11569_), .B(_11563_), .C(_11567_), .Y(_11576_) );
NAND3X1 NAND3X1_2653 ( .gnd(gnd), .vdd(vdd), .A(_11236_), .B(_11574_), .C(_11576_), .Y(_11577_) );
AOI21X1 AOI21X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_11573_), .B(_11577_), .C(_11441_), .Y(_11578_) );
NAND3X1 NAND3X1_2654 ( .gnd(gnd), .vdd(vdd), .A(_11240_), .B(_11574_), .C(_11576_), .Y(_11579_) );
NAND3X1 NAND3X1_2655 ( .gnd(gnd), .vdd(vdd), .A(_11236_), .B(_11568_), .C(_11572_), .Y(_11580_) );
AOI21X1 AOI21X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_11579_), .B(_11580_), .C(_11440_), .Y(_11581_) );
OAI21X1 OAI21X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_11578_), .B(_11581_), .C(_9845_), .Y(_11582_) );
INVX1 INVX1_1570 ( .gnd(gnd), .vdd(vdd), .A(_9845_), .Y(_11583_) );
NAND3X1 NAND3X1_2656 ( .gnd(gnd), .vdd(vdd), .A(_11440_), .B(_11579_), .C(_11580_), .Y(_11584_) );
NAND3X1 NAND3X1_2657 ( .gnd(gnd), .vdd(vdd), .A(_11573_), .B(_11577_), .C(_11441_), .Y(_11585_) );
NAND3X1 NAND3X1_2658 ( .gnd(gnd), .vdd(vdd), .A(_11583_), .B(_11584_), .C(_11585_), .Y(_11587_) );
NAND3X1 NAND3X1_2659 ( .gnd(gnd), .vdd(vdd), .A(_9884_), .B(_11587_), .C(_11582_), .Y(_11588_) );
NAND2X1 NAND2X1_1478 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_142_), .B(_11588_), .Y(_11589_) );
INVX1 INVX1_1571 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_142_), .Y(_11590_) );
OAI21X1 OAI21X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_11578_), .B(_11581_), .C(_11583_), .Y(_11591_) );
NAND3X1 NAND3X1_2660 ( .gnd(gnd), .vdd(vdd), .A(_9845_), .B(_11584_), .C(_11585_), .Y(_11592_) );
NAND2X1 NAND2X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_11592_), .B(_11591_), .Y(_11593_) );
NAND3X1 NAND3X1_2661 ( .gnd(gnd), .vdd(vdd), .A(_11590_), .B(_9884_), .C(_11593_), .Y(_11594_) );
NAND3X1 NAND3X1_2662 ( .gnd(gnd), .vdd(vdd), .A(_11253_), .B(_11594_), .C(_11589_), .Y(_11595_) );
INVX1 INVX1_1572 ( .gnd(gnd), .vdd(vdd), .A(_11253_), .Y(_11596_) );
NAND3X1 NAND3X1_2663 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_142_), .B(_9884_), .C(_11593_), .Y(_11598_) );
NAND2X1 NAND2X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_11590_), .B(_11588_), .Y(_11599_) );
NAND3X1 NAND3X1_2664 ( .gnd(gnd), .vdd(vdd), .A(_11596_), .B(_11598_), .C(_11599_), .Y(_11600_) );
NAND3X1 NAND3X1_2665 ( .gnd(gnd), .vdd(vdd), .A(_11439_), .B(_11595_), .C(_11600_), .Y(_11601_) );
INVX1 INVX1_1573 ( .gnd(gnd), .vdd(vdd), .A(_11439_), .Y(_11602_) );
NAND3X1 NAND3X1_2666 ( .gnd(gnd), .vdd(vdd), .A(_11596_), .B(_11594_), .C(_11589_), .Y(_11603_) );
NAND3X1 NAND3X1_2667 ( .gnd(gnd), .vdd(vdd), .A(_11253_), .B(_11598_), .C(_11599_), .Y(_11604_) );
NAND3X1 NAND3X1_2668 ( .gnd(gnd), .vdd(vdd), .A(_11602_), .B(_11603_), .C(_11604_), .Y(_11605_) );
NAND3X1 NAND3X1_2669 ( .gnd(gnd), .vdd(vdd), .A(_9572_), .B(_11601_), .C(_11605_), .Y(_11606_) );
AOI21X1 AOI21X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_11603_), .B(_11604_), .C(_11602_), .Y(_11607_) );
AOI21X1 AOI21X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_11595_), .B(_11600_), .C(_11439_), .Y(_11609_) );
OAI21X1 OAI21X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_11607_), .B(_11609_), .C(_9571_), .Y(_11610_) );
NAND3X1 NAND3X1_2670 ( .gnd(gnd), .vdd(vdd), .A(_9918_), .B(_11606_), .C(_11610_), .Y(_11611_) );
NAND2X1 NAND2X1_1481 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_158_), .B(_11611_), .Y(_11612_) );
INVX1 INVX1_1574 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_158_), .Y(_11613_) );
NAND2X1 NAND2X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_11601_), .B(_11605_), .Y(_11614_) );
AOI21X1 AOI21X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_9571_), .B(_11614_), .C(_9919_), .Y(_11615_) );
NAND3X1 NAND3X1_2671 ( .gnd(gnd), .vdd(vdd), .A(_11613_), .B(_11606_), .C(_11615_), .Y(_11616_) );
NAND3X1 NAND3X1_2672 ( .gnd(gnd), .vdd(vdd), .A(_11438_), .B(_11616_), .C(_11612_), .Y(_11617_) );
NAND3X1 NAND3X1_2673 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_158_), .B(_11606_), .C(_11615_), .Y(_11618_) );
NAND2X1 NAND2X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_11613_), .B(_11611_), .Y(_11620_) );
NAND3X1 NAND3X1_2674 ( .gnd(gnd), .vdd(vdd), .A(_11275_), .B(_11618_), .C(_11620_), .Y(_11621_) );
AOI21X1 AOI21X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_11617_), .B(_11621_), .C(_11437_), .Y(_11622_) );
NAND3X1 NAND3X1_2675 ( .gnd(gnd), .vdd(vdd), .A(_11275_), .B(_11616_), .C(_11612_), .Y(_11623_) );
NAND3X1 NAND3X1_2676 ( .gnd(gnd), .vdd(vdd), .A(_11438_), .B(_11618_), .C(_11620_), .Y(_11624_) );
AOI21X1 AOI21X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_11623_), .B(_11624_), .C(_11436_), .Y(_11625_) );
OAI21X1 OAI21X1_1841 ( .gnd(gnd), .vdd(vdd), .A(_11622_), .B(_11625_), .C(_12184_), .Y(_11626_) );
NAND3X1 NAND3X1_2677 ( .gnd(gnd), .vdd(vdd), .A(_11436_), .B(_11623_), .C(_11624_), .Y(_11627_) );
NAND3X1 NAND3X1_2678 ( .gnd(gnd), .vdd(vdd), .A(_11437_), .B(_11617_), .C(_11621_), .Y(_11628_) );
NAND3X1 NAND3X1_2679 ( .gnd(gnd), .vdd(vdd), .A(_12397_), .B(_11627_), .C(_11628_), .Y(_11629_) );
NAND3X1 NAND3X1_2680 ( .gnd(gnd), .vdd(vdd), .A(_9953_), .B(_11629_), .C(_11626_), .Y(_11631_) );
NAND2X1 NAND2X1_1484 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_174_), .B(_11631_), .Y(_11632_) );
INVX1 INVX1_1575 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_174_), .Y(_11633_) );
OAI21X1 OAI21X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_11622_), .B(_11625_), .C(_12397_), .Y(_11634_) );
NAND3X1 NAND3X1_2681 ( .gnd(gnd), .vdd(vdd), .A(_12184_), .B(_11627_), .C(_11628_), .Y(_11635_) );
NAND2X1 NAND2X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_11635_), .B(_11634_), .Y(_11636_) );
NAND3X1 NAND3X1_2682 ( .gnd(gnd), .vdd(vdd), .A(_11633_), .B(_9953_), .C(_11636_), .Y(_11637_) );
NAND3X1 NAND3X1_2683 ( .gnd(gnd), .vdd(vdd), .A(_11435_), .B(_11637_), .C(_11632_), .Y(_11638_) );
NAND3X1 NAND3X1_2684 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_174_), .B(_9953_), .C(_11636_), .Y(_11639_) );
NAND2X1 NAND2X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_11633_), .B(_11631_), .Y(_11640_) );
NAND3X1 NAND3X1_2685 ( .gnd(gnd), .vdd(vdd), .A(_11297_), .B(_11639_), .C(_11640_), .Y(_11642_) );
AOI21X1 AOI21X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_11638_), .B(_11642_), .C(_11434_), .Y(_11643_) );
NAND3X1 NAND3X1_2686 ( .gnd(gnd), .vdd(vdd), .A(_11297_), .B(_11637_), .C(_11632_), .Y(_11644_) );
NAND3X1 NAND3X1_2687 ( .gnd(gnd), .vdd(vdd), .A(_11435_), .B(_11639_), .C(_11640_), .Y(_11645_) );
AOI21X1 AOI21X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_11644_), .B(_11645_), .C(_11433_), .Y(_11646_) );
OAI21X1 OAI21X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_11646_), .B(_11643_), .C(_12194_), .Y(_11647_) );
NAND3X1 NAND3X1_2688 ( .gnd(gnd), .vdd(vdd), .A(_11433_), .B(_11644_), .C(_11645_), .Y(_11648_) );
NAND3X1 NAND3X1_2689 ( .gnd(gnd), .vdd(vdd), .A(_11638_), .B(_11434_), .C(_11642_), .Y(_11649_) );
NAND3X1 NAND3X1_2690 ( .gnd(gnd), .vdd(vdd), .A(_9566_), .B(_11648_), .C(_11649_), .Y(_11650_) );
NAND3X1 NAND3X1_2691 ( .gnd(gnd), .vdd(vdd), .A(_9991_), .B(_11650_), .C(_11647_), .Y(_11651_) );
NAND2X1 NAND2X1_1487 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_190_), .B(_11651_), .Y(_11653_) );
INVX1 INVX1_1576 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_190_), .Y(_11654_) );
OAI21X1 OAI21X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_11646_), .B(_11643_), .C(_9566_), .Y(_11655_) );
NAND3X1 NAND3X1_2692 ( .gnd(gnd), .vdd(vdd), .A(_12194_), .B(_11648_), .C(_11649_), .Y(_11656_) );
NAND2X1 NAND2X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_11656_), .B(_11655_), .Y(_11657_) );
NAND3X1 NAND3X1_2693 ( .gnd(gnd), .vdd(vdd), .A(_11654_), .B(_9991_), .C(_11657_), .Y(_11658_) );
NAND3X1 NAND3X1_2694 ( .gnd(gnd), .vdd(vdd), .A(_11431_), .B(_11658_), .C(_11653_), .Y(_11659_) );
NAND3X1 NAND3X1_2695 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_190_), .B(_9991_), .C(_11657_), .Y(_11660_) );
NAND2X1 NAND2X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_11654_), .B(_11651_), .Y(_11661_) );
NAND3X1 NAND3X1_2696 ( .gnd(gnd), .vdd(vdd), .A(_11327_), .B(_11660_), .C(_11661_), .Y(_11662_) );
AOI21X1 AOI21X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_11659_), .B(_11662_), .C(_11430_), .Y(_11664_) );
NAND3X1 NAND3X1_2697 ( .gnd(gnd), .vdd(vdd), .A(_11327_), .B(_11658_), .C(_11653_), .Y(_11665_) );
NAND3X1 NAND3X1_2698 ( .gnd(gnd), .vdd(vdd), .A(_11431_), .B(_11660_), .C(_11661_), .Y(_11666_) );
AOI21X1 AOI21X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_11665_), .B(_11666_), .C(_11429_), .Y(_11667_) );
OAI21X1 OAI21X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_11664_), .B(_11667_), .C(_9562_), .Y(_11668_) );
NAND3X1 NAND3X1_2699 ( .gnd(gnd), .vdd(vdd), .A(_11429_), .B(_11665_), .C(_11666_), .Y(_11669_) );
NAND3X1 NAND3X1_2700 ( .gnd(gnd), .vdd(vdd), .A(_11659_), .B(_11662_), .C(_11430_), .Y(_11670_) );
NAND3X1 NAND3X1_2701 ( .gnd(gnd), .vdd(vdd), .A(_9563_), .B(_11669_), .C(_11670_), .Y(_11671_) );
NAND3X1 NAND3X1_2702 ( .gnd(gnd), .vdd(vdd), .A(_10027_), .B(_11671_), .C(_11668_), .Y(_11672_) );
NAND2X1 NAND2X1_1490 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_206_), .B(_11672_), .Y(_11673_) );
INVX1 INVX1_1577 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_206_), .Y(_11675_) );
NAND3X1 NAND3X1_2703 ( .gnd(gnd), .vdd(vdd), .A(_9562_), .B(_11669_), .C(_11670_), .Y(_11676_) );
OAI21X1 OAI21X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_11664_), .B(_11667_), .C(_9563_), .Y(_11677_) );
NAND2X1 NAND2X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_11676_), .B(_11677_), .Y(_11678_) );
NAND3X1 NAND3X1_2704 ( .gnd(gnd), .vdd(vdd), .A(_11675_), .B(_10027_), .C(_11678_), .Y(_11679_) );
NAND3X1 NAND3X1_2705 ( .gnd(gnd), .vdd(vdd), .A(_11342_), .B(_11679_), .C(_11673_), .Y(_11680_) );
INVX1 INVX1_1578 ( .gnd(gnd), .vdd(vdd), .A(_11342_), .Y(_11681_) );
NAND3X1 NAND3X1_2706 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_206_), .B(_10027_), .C(_11678_), .Y(_11682_) );
NAND2X1 NAND2X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_11675_), .B(_11672_), .Y(_11683_) );
NAND3X1 NAND3X1_2707 ( .gnd(gnd), .vdd(vdd), .A(_11681_), .B(_11682_), .C(_11683_), .Y(_11684_) );
NAND3X1 NAND3X1_2708 ( .gnd(gnd), .vdd(vdd), .A(_11428_), .B(_11680_), .C(_11684_), .Y(_11686_) );
AOI21X1 AOI21X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_11357_), .B(_11354_), .C(_11348_), .Y(_11687_) );
AOI21X1 AOI21X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_11682_), .B(_11683_), .C(_11681_), .Y(_11688_) );
AOI21X1 AOI21X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_11679_), .B(_11673_), .C(_11342_), .Y(_11689_) );
OAI21X1 OAI21X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_11688_), .B(_11689_), .C(_11687_), .Y(_11690_) );
NAND3X1 NAND3X1_2709 ( .gnd(gnd), .vdd(vdd), .A(_9559_), .B(_11686_), .C(_11690_), .Y(_11691_) );
NOR3X1 NOR3X1_336 ( .gnd(gnd), .vdd(vdd), .A(_11688_), .B(_11687_), .C(_11689_), .Y(_11692_) );
AOI21X1 AOI21X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_11680_), .B(_11684_), .C(_11428_), .Y(_11693_) );
OAI21X1 OAI21X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_11692_), .B(_11693_), .C(_12212_), .Y(_11694_) );
NAND3X1 NAND3X1_2710 ( .gnd(gnd), .vdd(vdd), .A(_10064_), .B(_11691_), .C(_11694_), .Y(_11695_) );
NAND2X1 NAND2X1_1493 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_222_), .B(_11695_), .Y(_11697_) );
INVX1 INVX1_1579 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_222_), .Y(_11698_) );
NAND2X1 NAND2X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_11686_), .B(_11690_), .Y(_11699_) );
AOI21X1 AOI21X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_12212_), .B(_11699_), .C(_10065_), .Y(_11700_) );
NAND3X1 NAND3X1_2711 ( .gnd(gnd), .vdd(vdd), .A(_11698_), .B(_11691_), .C(_11700_), .Y(_11701_) );
NAND3X1 NAND3X1_2712 ( .gnd(gnd), .vdd(vdd), .A(_11371_), .B(_11701_), .C(_11697_), .Y(_11702_) );
INVX1 INVX1_1580 ( .gnd(gnd), .vdd(vdd), .A(_11371_), .Y(_11703_) );
NAND3X1 NAND3X1_2713 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_222_), .B(_11691_), .C(_11700_), .Y(_11704_) );
NAND2X1 NAND2X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_11698_), .B(_11695_), .Y(_11705_) );
NAND3X1 NAND3X1_2714 ( .gnd(gnd), .vdd(vdd), .A(_11703_), .B(_11704_), .C(_11705_), .Y(_11706_) );
NAND3X1 NAND3X1_2715 ( .gnd(gnd), .vdd(vdd), .A(_11427_), .B(_11702_), .C(_11706_), .Y(_11708_) );
AOI21X1 AOI21X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_11373_), .B(_11062_), .C(_11376_), .Y(_11709_) );
NAND3X1 NAND3X1_2716 ( .gnd(gnd), .vdd(vdd), .A(_11703_), .B(_11701_), .C(_11697_), .Y(_11710_) );
NAND3X1 NAND3X1_2717 ( .gnd(gnd), .vdd(vdd), .A(_11371_), .B(_11704_), .C(_11705_), .Y(_11711_) );
NAND3X1 NAND3X1_2718 ( .gnd(gnd), .vdd(vdd), .A(_11709_), .B(_11710_), .C(_11711_), .Y(_11712_) );
NAND3X1 NAND3X1_2719 ( .gnd(gnd), .vdd(vdd), .A(_9556_), .B(_11708_), .C(_11712_), .Y(_11713_) );
AOI21X1 AOI21X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_11710_), .B(_11711_), .C(_11709_), .Y(_11714_) );
AOI21X1 AOI21X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_11702_), .B(_11706_), .C(_11427_), .Y(_11715_) );
OAI21X1 OAI21X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_11714_), .B(_11715_), .C(_9555_), .Y(_11716_) );
NAND3X1 NAND3X1_2720 ( .gnd(gnd), .vdd(vdd), .A(_10101_), .B(_11713_), .C(_11716_), .Y(_11717_) );
NAND2X1 NAND2X1_1496 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_238_), .B(_11717_), .Y(_11719_) );
INVX1 INVX1_1581 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_238_), .Y(_11720_) );
NAND2X1 NAND2X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_11708_), .B(_11712_), .Y(_11721_) );
AOI21X1 AOI21X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_9555_), .B(_11721_), .C(_10102_), .Y(_11722_) );
NAND3X1 NAND3X1_2721 ( .gnd(gnd), .vdd(vdd), .A(_11720_), .B(_11713_), .C(_11722_), .Y(_11723_) );
NAND3X1 NAND3X1_2722 ( .gnd(gnd), .vdd(vdd), .A(_11386_), .B(_11723_), .C(_11719_), .Y(_11724_) );
INVX2 INVX2_381 ( .gnd(gnd), .vdd(vdd), .A(_11386_), .Y(_11725_) );
NAND3X1 NAND3X1_2723 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_238_), .B(_11713_), .C(_11722_), .Y(_11726_) );
NAND2X1 NAND2X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_11720_), .B(_11717_), .Y(_11727_) );
NAND3X1 NAND3X1_2724 ( .gnd(gnd), .vdd(vdd), .A(_11725_), .B(_11726_), .C(_11727_), .Y(_11728_) );
NAND3X1 NAND3X1_2725 ( .gnd(gnd), .vdd(vdd), .A(_11724_), .B(_11728_), .C(_11426_), .Y(_11730_) );
AOI21X1 AOI21X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_11401_), .B(_11398_), .C(_11392_), .Y(_11731_) );
AOI21X1 AOI21X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_11726_), .B(_11727_), .C(_11725_), .Y(_11732_) );
AOI21X1 AOI21X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_11723_), .B(_11719_), .C(_11386_), .Y(_11733_) );
OAI21X1 OAI21X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_11732_), .B(_11733_), .C(_11731_), .Y(_11734_) );
NAND3X1 NAND3X1_2726 ( .gnd(gnd), .vdd(vdd), .A(_12462_), .B(_11730_), .C(_11734_), .Y(_11735_) );
NAND3X1 NAND3X1_2727 ( .gnd(gnd), .vdd(vdd), .A(_11725_), .B(_11723_), .C(_11719_), .Y(_11736_) );
NAND3X1 NAND3X1_2728 ( .gnd(gnd), .vdd(vdd), .A(_11386_), .B(_11726_), .C(_11727_), .Y(_11737_) );
AOI21X1 AOI21X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_11736_), .B(_11737_), .C(_11731_), .Y(_11738_) );
AOI21X1 AOI21X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_11724_), .B(_11728_), .C(_11426_), .Y(_11739_) );
OAI21X1 OAI21X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_11738_), .B(_11739_), .C(_12234_), .Y(_11741_) );
NAND3X1 NAND3X1_2729 ( .gnd(gnd), .vdd(vdd), .A(_10136_), .B(_11735_), .C(_11741_), .Y(_11742_) );
NAND2X1 NAND2X1_1499 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_254_), .B(_11742_), .Y(_11743_) );
INVX1 INVX1_1582 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_254_), .Y(_11744_) );
NAND2X1 NAND2X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_11730_), .B(_11734_), .Y(_11745_) );
AOI21X1 AOI21X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_12234_), .B(_11745_), .C(_10137_), .Y(_11746_) );
NAND3X1 NAND3X1_2730 ( .gnd(gnd), .vdd(vdd), .A(_11744_), .B(_11735_), .C(_11746_), .Y(_11747_) );
NAND3X1 NAND3X1_2731 ( .gnd(gnd), .vdd(vdd), .A(_11425_), .B(_11747_), .C(_11743_), .Y(_11748_) );
INVX1 INVX1_1583 ( .gnd(gnd), .vdd(vdd), .A(_11748_), .Y(_11749_) );
AOI21X1 AOI21X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_11747_), .B(_11743_), .C(_11425_), .Y(_11750_) );
OAI21X1 OAI21X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_11749_), .B(_11750_), .C(_11424_), .Y(_11752_) );
INVX1 INVX1_1584 ( .gnd(gnd), .vdd(vdd), .A(_11750_), .Y(_11753_) );
NAND3X1 NAND3X1_2732 ( .gnd(gnd), .vdd(vdd), .A(_11423_), .B(_11748_), .C(_11753_), .Y(_11754_) );
NAND2X1 NAND2X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_11752_), .B(_11754_), .Y(module_2_H_22_) );
OAI21X1 OAI21X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_11423_), .B(_11750_), .C(_11748_), .Y(_11755_) );
AOI21X1 AOI21X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_11735_), .B(_11746_), .C(_11744_), .Y(_11756_) );
INVX1 INVX1_1585 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_255_), .Y(_11757_) );
OAI21X1 OAI21X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_11731_), .B(_11733_), .C(_11724_), .Y(_11758_) );
INVX1 INVX1_1586 ( .gnd(gnd), .vdd(vdd), .A(_11758_), .Y(_11759_) );
NAND2X1 NAND2X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_11702_), .B(_11708_), .Y(_11760_) );
OAI21X1 OAI21X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_11689_), .B(_11687_), .C(_11680_), .Y(_11762_) );
NAND2X1 NAND2X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_11665_), .B(_11669_), .Y(_11763_) );
NAND2X1 NAND2X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_11644_), .B(_11648_), .Y(_11764_) );
INVX1 INVX1_1587 ( .gnd(gnd), .vdd(vdd), .A(_11764_), .Y(_11765_) );
NAND2X1 NAND2X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_11623_), .B(_11627_), .Y(_11766_) );
NAND2X1 NAND2X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_11595_), .B(_11601_), .Y(_11767_) );
NAND2X1 NAND2X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_11579_), .B(_11584_), .Y(_11768_) );
INVX1 INVX1_1588 ( .gnd(gnd), .vdd(vdd), .A(_11768_), .Y(_11769_) );
INVX1 INVX1_1589 ( .gnd(gnd), .vdd(vdd), .A(_11574_), .Y(_11770_) );
NOR2X1 NOR2X1_853 ( .gnd(gnd), .vdd(vdd), .A(_12368_), .B(_12370_), .Y(_11771_) );
NAND2X1 NAND2X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_11551_), .B(_11556_), .Y(_11773_) );
INVX1 INVX1_1590 ( .gnd(gnd), .vdd(vdd), .A(_11773_), .Y(_11774_) );
OAI21X1 OAI21X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_11537_), .B(_11535_), .C(_11529_), .Y(_11775_) );
INVX1 INVX1_1591 ( .gnd(gnd), .vdd(vdd), .A(_12350_), .Y(_11776_) );
NAND2X1 NAND2X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_11507_), .B(_11512_), .Y(_11777_) );
INVX1 INVX1_1592 ( .gnd(gnd), .vdd(vdd), .A(_11777_), .Y(_11778_) );
NAND2X1 NAND2X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_11485_), .B(_11490_), .Y(_11779_) );
INVX1 INVX1_1593 ( .gnd(gnd), .vdd(vdd), .A(_10388_), .Y(_11780_) );
XNOR2X1 XNOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_11480_), .B(_11780_), .Y(_11781_) );
INVX1 INVX1_1594 ( .gnd(gnd), .vdd(vdd), .A(_11781_), .Y(_11782_) );
INVX1 INVX1_1595 ( .gnd(gnd), .vdd(vdd), .A(_11447_), .Y(_11784_) );
NAND2X1 NAND2X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_11467_), .B(_11470_), .Y(_11785_) );
OAI21X1 OAI21X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_11785_), .B(_11784_), .C(_11467_), .Y(_11786_) );
INVX1 INVX1_1596 ( .gnd(gnd), .vdd(vdd), .A(_11786_), .Y(_11787_) );
INVX1 INVX1_1597 ( .gnd(gnd), .vdd(vdd), .A(_11462_), .Y(_11788_) );
OAI21X1 OAI21X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_11118_), .B(_11123_), .C(_11458_), .Y(_11789_) );
OAI21X1 OAI21X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_11112_), .B(_11457_), .C(_11789_), .Y(_11790_) );
INVX1 INVX1_1598 ( .gnd(gnd), .vdd(vdd), .A(_11790_), .Y(_11791_) );
OAI21X1 OAI21X1_1860 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_12_), .B(module_2_W_13_), .C(module_2_W_14_), .Y(_11792_) );
XOR2X1 XOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_11_), .B(module_2_W_15_), .Y(_11793_) );
XNOR2X1 XNOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_11793_), .B(_11792_), .Y(_11795_) );
XOR2X1 XOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_12285_), .B(module_2_W_31_), .Y(_11796_) );
XNOR2X1 XNOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_11796_), .B(_11795_), .Y(_11797_) );
XOR2X1 XOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_11455_), .B(_11797_), .Y(_11798_) );
XNOR2X1 XNOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_11798_), .B(_10184_), .Y(_11799_) );
XNOR2X1 XNOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_10352_), .B(bloque_datos[15]), .Y(_11800_) );
XNOR2X1 XNOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_11799_), .B(_11800_), .Y(_11801_) );
NOR2X1 NOR2X1_854 ( .gnd(gnd), .vdd(vdd), .A(_11791_), .B(_11801_), .Y(_11802_) );
NAND2X1 NAND2X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_11791_), .B(_11801_), .Y(_11803_) );
INVX1 INVX1_1599 ( .gnd(gnd), .vdd(vdd), .A(_11803_), .Y(_11804_) );
OR2X2 OR2X2_256 ( .gnd(gnd), .vdd(vdd), .A(_11804_), .B(_11802_), .Y(_11806_) );
NOR2X1 NOR2X1_855 ( .gnd(gnd), .vdd(vdd), .A(_11788_), .B(_11806_), .Y(_11807_) );
INVX1 INVX1_1600 ( .gnd(gnd), .vdd(vdd), .A(_11807_), .Y(_11808_) );
OAI21X1 OAI21X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_11804_), .B(_11802_), .C(_11788_), .Y(_11809_) );
XNOR2X1 XNOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_10366_), .B(_10190_), .Y(_11810_) );
INVX1 INVX1_1601 ( .gnd(gnd), .vdd(vdd), .A(_11810_), .Y(_11811_) );
NAND3X1 NAND3X1_2733 ( .gnd(gnd), .vdd(vdd), .A(_11809_), .B(_11811_), .C(_11808_), .Y(_11812_) );
AOI21X1 AOI21X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_11809_), .B(_11808_), .C(_11811_), .Y(_11813_) );
INVX1 INVX1_1602 ( .gnd(gnd), .vdd(vdd), .A(_11813_), .Y(_11814_) );
NAND2X1 NAND2X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_11812_), .B(_11814_), .Y(_11815_) );
NOR2X1 NOR2X1_856 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf3_), .B(_11815_), .Y(_11817_) );
AND2X2 AND2X2_247 ( .gnd(gnd), .vdd(vdd), .A(_11815_), .B(bloque_datos_31_bF_buf2_), .Y(_11818_) );
NOR2X1 NOR2X1_857 ( .gnd(gnd), .vdd(vdd), .A(_11817_), .B(_11818_), .Y(_11819_) );
NAND2X1 NAND2X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_11787_), .B(_11819_), .Y(_11820_) );
OAI21X1 OAI21X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_11818_), .B(_11817_), .C(_11786_), .Y(_11821_) );
XOR2X1 XOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_10205_), .B(bloque_datos_47_bF_buf3_), .Y(_11822_) );
NAND3X1 NAND3X1_2734 ( .gnd(gnd), .vdd(vdd), .A(_11821_), .B(_11822_), .C(_11820_), .Y(_11823_) );
AND2X2 AND2X2_248 ( .gnd(gnd), .vdd(vdd), .A(_11819_), .B(_11787_), .Y(_11824_) );
NOR2X1 NOR2X1_858 ( .gnd(gnd), .vdd(vdd), .A(_11787_), .B(_11819_), .Y(_11825_) );
INVX1 INVX1_1603 ( .gnd(gnd), .vdd(vdd), .A(_11822_), .Y(_11826_) );
OAI21X1 OAI21X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_11824_), .B(_11825_), .C(_11826_), .Y(_11828_) );
AOI21X1 AOI21X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_11823_), .B(_11828_), .C(_11782_), .Y(_11829_) );
INVX1 INVX1_1604 ( .gnd(gnd), .vdd(vdd), .A(_11829_), .Y(_11830_) );
NAND3X1 NAND3X1_2735 ( .gnd(gnd), .vdd(vdd), .A(_11782_), .B(_11823_), .C(_11828_), .Y(_11831_) );
NAND3X1 NAND3X1_2736 ( .gnd(gnd), .vdd(vdd), .A(_11779_), .B(_11831_), .C(_11830_), .Y(_11832_) );
INVX1 INVX1_1605 ( .gnd(gnd), .vdd(vdd), .A(_11779_), .Y(_11833_) );
INVX1 INVX1_1606 ( .gnd(gnd), .vdd(vdd), .A(_11831_), .Y(_11834_) );
OAI21X1 OAI21X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_11834_), .B(_11829_), .C(_11833_), .Y(_11835_) );
OAI21X1 OAI21X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_10216_), .B(_10213_), .C(_12506_), .Y(_11836_) );
NAND2X1 NAND2X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_12335_), .B(_10340_), .Y(_11837_) );
NAND2X1 NAND2X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_11836_), .B(_11837_), .Y(_11839_) );
AOI21X1 AOI21X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_11835_), .B(_11832_), .C(_11839_), .Y(_11840_) );
NAND3X1 NAND3X1_2737 ( .gnd(gnd), .vdd(vdd), .A(_11833_), .B(_11831_), .C(_11830_), .Y(_11841_) );
OAI21X1 OAI21X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_11834_), .B(_11829_), .C(_11779_), .Y(_11842_) );
AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_11836_), .B(_11837_), .C(_11841_), .D(_11842_), .Y(_11843_) );
NOR2X1 NOR2X1_859 ( .gnd(gnd), .vdd(vdd), .A(_11840_), .B(_11843_), .Y(_11844_) );
XNOR2X1 XNOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_11502_), .B(bloque_datos[63]), .Y(_11845_) );
AND2X2 AND2X2_249 ( .gnd(gnd), .vdd(vdd), .A(_11844_), .B(_11845_), .Y(_11846_) );
NOR2X1 NOR2X1_860 ( .gnd(gnd), .vdd(vdd), .A(_11845_), .B(_11844_), .Y(_11847_) );
OAI21X1 OAI21X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_11846_), .B(_11847_), .C(_11778_), .Y(_11848_) );
NAND2X1 NAND2X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_11845_), .B(_11844_), .Y(_11850_) );
OR2X2 OR2X2_257 ( .gnd(gnd), .vdd(vdd), .A(_11844_), .B(_11845_), .Y(_11851_) );
NAND3X1 NAND3X1_2738 ( .gnd(gnd), .vdd(vdd), .A(_11777_), .B(_11850_), .C(_11851_), .Y(_11852_) );
NAND3X1 NAND3X1_2739 ( .gnd(gnd), .vdd(vdd), .A(_11776_), .B(_11848_), .C(_11852_), .Y(_11853_) );
NAND3X1 NAND3X1_2740 ( .gnd(gnd), .vdd(vdd), .A(_11778_), .B(_11850_), .C(_11851_), .Y(_11854_) );
OAI21X1 OAI21X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_11846_), .B(_11847_), .C(_11777_), .Y(_11855_) );
NAND3X1 NAND3X1_2741 ( .gnd(gnd), .vdd(vdd), .A(_12350_), .B(_11855_), .C(_11854_), .Y(_11856_) );
NAND2X1 NAND2X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_11853_), .B(_11856_), .Y(_11857_) );
XOR2X1 XOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_10338_), .B(bloque_datos_79_bF_buf3_), .Y(_11858_) );
NOR2X1 NOR2X1_861 ( .gnd(gnd), .vdd(vdd), .A(_11524_), .B(_11858_), .Y(_11859_) );
INVX1 INVX1_1607 ( .gnd(gnd), .vdd(vdd), .A(_11859_), .Y(_11861_) );
NAND2X1 NAND2X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_11524_), .B(_11858_), .Y(_11862_) );
NAND2X1 NAND2X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_11862_), .B(_11861_), .Y(_11863_) );
NAND2X1 NAND2X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_11863_), .B(_11857_), .Y(_11864_) );
OR2X2 OR2X2_258 ( .gnd(gnd), .vdd(vdd), .A(_11857_), .B(_11863_), .Y(_11865_) );
NAND3X1 NAND3X1_2742 ( .gnd(gnd), .vdd(vdd), .A(_11775_), .B(_11864_), .C(_11865_), .Y(_11866_) );
INVX1 INVX1_1608 ( .gnd(gnd), .vdd(vdd), .A(_11775_), .Y(_11867_) );
AND2X2 AND2X2_250 ( .gnd(gnd), .vdd(vdd), .A(_11857_), .B(_11863_), .Y(_11868_) );
NOR2X1 NOR2X1_862 ( .gnd(gnd), .vdd(vdd), .A(_11863_), .B(_11857_), .Y(_11869_) );
OAI21X1 OAI21X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_11868_), .B(_11869_), .C(_11867_), .Y(_11870_) );
NOR2X1 NOR2X1_863 ( .gnd(gnd), .vdd(vdd), .A(_12356_), .B(_12358_), .Y(_11872_) );
XNOR2X1 XNOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_10336_), .B(_11872_), .Y(_11873_) );
INVX1 INVX1_1609 ( .gnd(gnd), .vdd(vdd), .A(_11873_), .Y(_11874_) );
AOI21X1 AOI21X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_11870_), .B(_11866_), .C(_11874_), .Y(_11875_) );
NAND3X1 NAND3X1_2743 ( .gnd(gnd), .vdd(vdd), .A(_11867_), .B(_11864_), .C(_11865_), .Y(_11876_) );
OAI21X1 OAI21X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_11868_), .B(_11869_), .C(_11775_), .Y(_11877_) );
AOI21X1 AOI21X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_11877_), .B(_11876_), .C(_11873_), .Y(_11878_) );
NOR2X1 NOR2X1_864 ( .gnd(gnd), .vdd(vdd), .A(_11875_), .B(_11878_), .Y(_11879_) );
NAND2X1 NAND2X1_1522 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf3_), .B(_11546_), .Y(_11880_) );
NOR2X1 NOR2X1_865 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf2_), .B(_11546_), .Y(_11881_) );
INVX1 INVX1_1610 ( .gnd(gnd), .vdd(vdd), .A(_11881_), .Y(_11883_) );
NAND2X1 NAND2X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_11880_), .B(_11883_), .Y(_11884_) );
NAND2X1 NAND2X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_11884_), .B(_11879_), .Y(_11885_) );
OR2X2 OR2X2_259 ( .gnd(gnd), .vdd(vdd), .A(_11879_), .B(_11884_), .Y(_11886_) );
NAND3X1 NAND3X1_2744 ( .gnd(gnd), .vdd(vdd), .A(_11774_), .B(_11885_), .C(_11886_), .Y(_11887_) );
AND2X2 AND2X2_251 ( .gnd(gnd), .vdd(vdd), .A(_11879_), .B(_11884_), .Y(_11888_) );
NOR2X1 NOR2X1_866 ( .gnd(gnd), .vdd(vdd), .A(_11884_), .B(_11879_), .Y(_11889_) );
OAI21X1 OAI21X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_11888_), .B(_11889_), .C(_11773_), .Y(_11890_) );
AOI21X1 AOI21X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_11890_), .B(_11887_), .C(_11771_), .Y(_11891_) );
INVX1 INVX1_1611 ( .gnd(gnd), .vdd(vdd), .A(_11771_), .Y(_11892_) );
OAI21X1 OAI21X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_11888_), .B(_11889_), .C(_11774_), .Y(_11894_) );
NAND3X1 NAND3X1_2745 ( .gnd(gnd), .vdd(vdd), .A(_11773_), .B(_11885_), .C(_11886_), .Y(_11895_) );
AOI21X1 AOI21X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_11894_), .B(_11895_), .C(_11892_), .Y(_11896_) );
OAI21X1 OAI21X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_11891_), .B(_11896_), .C(_11770_), .Y(_11897_) );
NAND3X1 NAND3X1_2746 ( .gnd(gnd), .vdd(vdd), .A(_11892_), .B(_11894_), .C(_11895_), .Y(_11898_) );
NAND3X1 NAND3X1_2747 ( .gnd(gnd), .vdd(vdd), .A(_11771_), .B(_11890_), .C(_11887_), .Y(_11899_) );
NAND3X1 NAND3X1_2748 ( .gnd(gnd), .vdd(vdd), .A(_11574_), .B(_11898_), .C(_11899_), .Y(_11900_) );
NAND2X1 NAND2X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_11900_), .B(_11897_), .Y(_11901_) );
AOI21X1 AOI21X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_11769_), .B(_11901_), .C(_10249_), .Y(_11902_) );
OAI21X1 OAI21X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_11769_), .B(_11901_), .C(_11902_), .Y(_11903_) );
XOR2X1 XOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_10505_), .B(module_2_W_143_), .Y(_11905_) );
XOR2X1 XOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_11903_), .B(_11905_), .Y(_11906_) );
XOR2X1 XOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_11906_), .B(_11589_), .Y(_11907_) );
NAND2X1 NAND2X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_11767_), .B(_11907_), .Y(_11908_) );
INVX1 INVX1_1612 ( .gnd(gnd), .vdd(vdd), .A(_11767_), .Y(_11909_) );
XNOR2X1 XNOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_11906_), .B(_11589_), .Y(_11910_) );
AOI21X1 AOI21X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_11909_), .B(_11910_), .C(_10503_), .Y(_11911_) );
XNOR2X1 XNOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_12393_), .B(module_2_W_159_), .Y(_11912_) );
NAND3X1 NAND3X1_2749 ( .gnd(gnd), .vdd(vdd), .A(_11908_), .B(_11912_), .C(_11911_), .Y(_11913_) );
NOR2X1 NOR2X1_867 ( .gnd(gnd), .vdd(vdd), .A(_11909_), .B(_11910_), .Y(_11914_) );
OAI21X1 OAI21X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_11907_), .B(_11767_), .C(_10258_), .Y(_11916_) );
INVX1 INVX1_1613 ( .gnd(gnd), .vdd(vdd), .A(_11912_), .Y(_11917_) );
OAI21X1 OAI21X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_11916_), .B(_11914_), .C(_11917_), .Y(_11918_) );
NAND2X1 NAND2X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_11913_), .B(_11918_), .Y(_11919_) );
XOR2X1 XOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_11919_), .B(_11612_), .Y(_11920_) );
NAND2X1 NAND2X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_11766_), .B(_11920_), .Y(_11921_) );
INVX1 INVX1_1614 ( .gnd(gnd), .vdd(vdd), .A(_11766_), .Y(_11922_) );
XNOR2X1 XNOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_11919_), .B(_11612_), .Y(_11923_) );
AOI21X1 AOI21X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_11922_), .B(_11923_), .C(_10271_), .Y(_11924_) );
XOR2X1 XOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_12404_), .B(module_2_W_175_), .Y(_11925_) );
NAND3X1 NAND3X1_2750 ( .gnd(gnd), .vdd(vdd), .A(_11921_), .B(_11925_), .C(_11924_), .Y(_11927_) );
NOR2X1 NOR2X1_868 ( .gnd(gnd), .vdd(vdd), .A(_11922_), .B(_11923_), .Y(_11928_) );
OAI21X1 OAI21X1_1877 ( .gnd(gnd), .vdd(vdd), .A(_11920_), .B(_11766_), .C(_10332_), .Y(_11929_) );
INVX1 INVX1_1615 ( .gnd(gnd), .vdd(vdd), .A(_11925_), .Y(_11930_) );
OAI21X1 OAI21X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_11929_), .B(_11928_), .C(_11930_), .Y(_11931_) );
NAND2X1 NAND2X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_11927_), .B(_11931_), .Y(_11932_) );
XNOR2X1 XNOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_11932_), .B(_11632_), .Y(_11933_) );
NAND2X1 NAND2X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_11765_), .B(_11933_), .Y(_11934_) );
XOR2X1 XOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_11932_), .B(_11632_), .Y(_11935_) );
AOI21X1 AOI21X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_11764_), .B(_11935_), .C(_10281_), .Y(_11936_) );
AND2X2 AND2X2_252 ( .gnd(gnd), .vdd(vdd), .A(_8986_), .B(module_2_W_191_), .Y(_11938_) );
NOR2X1 NOR2X1_869 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_191_), .B(_8986_), .Y(_11939_) );
NOR2X1 NOR2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_11939_), .B(_11938_), .Y(_11940_) );
NAND3X1 NAND3X1_2751 ( .gnd(gnd), .vdd(vdd), .A(_11934_), .B(_11940_), .C(_11936_), .Y(_11941_) );
NOR2X1 NOR2X1_871 ( .gnd(gnd), .vdd(vdd), .A(_11764_), .B(_11935_), .Y(_11942_) );
OAI21X1 OAI21X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_11933_), .B(_11765_), .C(_10328_), .Y(_11943_) );
OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_11938_), .B(_11939_), .C(_11943_), .D(_11942_), .Y(_11944_) );
NAND2X1 NAND2X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_11941_), .B(_11944_), .Y(_11945_) );
XOR2X1 XOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_11945_), .B(_11653_), .Y(_11946_) );
NAND2X1 NAND2X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_11763_), .B(_11946_), .Y(_11947_) );
INVX1 INVX1_1616 ( .gnd(gnd), .vdd(vdd), .A(_11763_), .Y(_11949_) );
XNOR2X1 XNOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_11945_), .B(_11653_), .Y(_11950_) );
AOI21X1 AOI21X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_11949_), .B(_11950_), .C(_10567_), .Y(_11951_) );
OAI21X1 OAI21X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_12425_), .B(_12428_), .C(module_2_W_207_), .Y(_11952_) );
INVX1 INVX1_1617 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_207_), .Y(_11953_) );
NAND3X1 NAND3X1_2752 ( .gnd(gnd), .vdd(vdd), .A(_11953_), .B(_12427_), .C(_12432_), .Y(_11954_) );
NAND2X1 NAND2X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_11954_), .B(_11952_), .Y(_11955_) );
INVX1 INVX1_1618 ( .gnd(gnd), .vdd(vdd), .A(_11955_), .Y(_11956_) );
NAND3X1 NAND3X1_2753 ( .gnd(gnd), .vdd(vdd), .A(_11947_), .B(_11956_), .C(_11951_), .Y(_11957_) );
NOR2X1 NOR2X1_872 ( .gnd(gnd), .vdd(vdd), .A(_11949_), .B(_11950_), .Y(_11958_) );
OAI21X1 OAI21X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_11946_), .B(_11763_), .C(_10290_), .Y(_11960_) );
OAI21X1 OAI21X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_11960_), .B(_11958_), .C(_11955_), .Y(_11961_) );
NAND2X1 NAND2X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_11957_), .B(_11961_), .Y(_11962_) );
XOR2X1 XOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_11962_), .B(_11673_), .Y(_11963_) );
XNOR2X1 XNOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_11963_), .B(_11762_), .Y(_11964_) );
OAI21X1 OAI21X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_12440_), .B(_12443_), .C(module_2_W_223_), .Y(_11965_) );
INVX1 INVX1_1619 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_223_), .Y(_11966_) );
NAND2X1 NAND2X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_11966_), .B(_12445_), .Y(_11967_) );
NAND2X1 NAND2X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_11965_), .B(_11967_), .Y(_11968_) );
NOR3X1 NOR3X1_337 ( .gnd(gnd), .vdd(vdd), .A(_11968_), .B(_10301_), .C(_11964_), .Y(_11969_) );
XOR2X1 XOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_11963_), .B(_11762_), .Y(_11971_) );
AND2X2 AND2X2_253 ( .gnd(gnd), .vdd(vdd), .A(_11967_), .B(_11965_), .Y(_11972_) );
AOI21X1 AOI21X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_10580_), .B(_11971_), .C(_11972_), .Y(_11973_) );
OAI21X1 OAI21X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_11969_), .B(_11973_), .C(_11697_), .Y(_11974_) );
INVX1 INVX1_1620 ( .gnd(gnd), .vdd(vdd), .A(_11697_), .Y(_11975_) );
NAND3X1 NAND3X1_2754 ( .gnd(gnd), .vdd(vdd), .A(_10580_), .B(_11971_), .C(_11972_), .Y(_11976_) );
OAI21X1 OAI21X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_11964_), .B(_10301_), .C(_11968_), .Y(_11977_) );
NAND3X1 NAND3X1_2755 ( .gnd(gnd), .vdd(vdd), .A(_11975_), .B(_11976_), .C(_11977_), .Y(_11978_) );
AND2X2 AND2X2_254 ( .gnd(gnd), .vdd(vdd), .A(_11974_), .B(_11978_), .Y(_11979_) );
NAND2X1 NAND2X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_11760_), .B(_11979_), .Y(_11980_) );
INVX1 INVX1_1621 ( .gnd(gnd), .vdd(vdd), .A(_11760_), .Y(_11982_) );
NAND2X1 NAND2X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_11978_), .B(_11974_), .Y(_11983_) );
AOI21X1 AOI21X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_11983_), .B(_11982_), .C(_10311_), .Y(_11984_) );
OAI21X1 OAI21X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_12456_), .B(_12451_), .C(module_2_W_239_), .Y(_11985_) );
INVX1 INVX1_1622 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_239_), .Y(_11986_) );
NAND3X1 NAND3X1_2756 ( .gnd(gnd), .vdd(vdd), .A(_11986_), .B(_12450_), .C(_12455_), .Y(_11987_) );
AND2X2 AND2X2_255 ( .gnd(gnd), .vdd(vdd), .A(_11985_), .B(_11987_), .Y(_11988_) );
NAND3X1 NAND3X1_2757 ( .gnd(gnd), .vdd(vdd), .A(_11980_), .B(_11984_), .C(_11988_), .Y(_11989_) );
NOR2X1 NOR2X1_873 ( .gnd(gnd), .vdd(vdd), .A(_11983_), .B(_11982_), .Y(_11990_) );
OAI21X1 OAI21X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_11979_), .B(_11760_), .C(_10324_), .Y(_11991_) );
NAND2X1 NAND2X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_11987_), .B(_11985_), .Y(_11993_) );
OAI21X1 OAI21X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_11991_), .B(_11990_), .C(_11993_), .Y(_11994_) );
NAND2X1 NAND2X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_11994_), .B(_11989_), .Y(_11995_) );
XNOR2X1 XNOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_11995_), .B(_11719_), .Y(_11996_) );
NOR2X1 NOR2X1_874 ( .gnd(gnd), .vdd(vdd), .A(_11759_), .B(_11996_), .Y(_11997_) );
XOR2X1 XOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_11995_), .B(_11719_), .Y(_11998_) );
OAI21X1 OAI21X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_11998_), .B(_11758_), .C(_10323_), .Y(_11999_) );
OAI21X1 OAI21X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_11999_), .B(_11997_), .C(_11757_), .Y(_12000_) );
OAI21X1 OAI21X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_11738_), .B(_11732_), .C(_11998_), .Y(_12001_) );
AOI21X1 AOI21X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_11759_), .B(_11996_), .C(_10322_), .Y(_12002_) );
NAND3X1 NAND3X1_2758 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_255_), .B(_12001_), .C(_12002_), .Y(_12004_) );
NAND3X1 NAND3X1_2759 ( .gnd(gnd), .vdd(vdd), .A(_11756_), .B(_12004_), .C(_12000_), .Y(_12005_) );
NAND3X1 NAND3X1_2760 ( .gnd(gnd), .vdd(vdd), .A(_11757_), .B(_12001_), .C(_12002_), .Y(_12006_) );
OAI21X1 OAI21X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_11999_), .B(_11997_), .C(module_2_W_255_), .Y(_12007_) );
NAND3X1 NAND3X1_2761 ( .gnd(gnd), .vdd(vdd), .A(_11743_), .B(_12006_), .C(_12007_), .Y(_12008_) );
NAND2X1 NAND2X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_12008_), .B(_12005_), .Y(_12009_) );
XNOR2X1 XNOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_11755_), .B(_12009_), .Y(module_2_H_23_) );
INVX1 INVX1_1623 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_241_), .Y(_10559_) );
AND2X2 AND2X2_256 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_0_), .B(module_2_W_16_), .Y(_10570_) );
NOR2X1 NOR2X1_875 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_0_), .B(module_2_W_16_), .Y(_10581_) );
OAI21X1 OAI21X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_10570_), .B(_10581_), .C(bloque_datos[0]), .Y(_10592_) );
INVX1 INVX1_1624 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(_10603_) );
NOR2X1 NOR2X1_876 ( .gnd(gnd), .vdd(vdd), .A(_10581_), .B(_10570_), .Y(_10614_) );
NAND2X1 NAND2X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_10603_), .B(_10614_), .Y(_10625_) );
NAND2X1 NAND2X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_10592_), .B(_10625_), .Y(_10636_) );
NAND2X1 NAND2X1_1544 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf3_), .B(_10636_), .Y(_10647_) );
OR2X2 OR2X2_260 ( .gnd(gnd), .vdd(vdd), .A(_10636_), .B(bloque_datos_16_bF_buf2_), .Y(_10658_) );
NAND2X1 NAND2X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_10647_), .B(_10658_), .Y(_10667_) );
NAND2X1 NAND2X1_1546 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf2_), .B(_10667_), .Y(_10676_) );
OR2X2 OR2X2_261 ( .gnd(gnd), .vdd(vdd), .A(_10667_), .B(bloque_datos_32_bF_buf1_), .Y(_10686_) );
NAND2X1 NAND2X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_10676_), .B(_10686_), .Y(_10697_) );
NAND2X1 NAND2X1_1548 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_48_bF_buf2_), .B(_10697_), .Y(_10708_) );
OR2X2 OR2X2_262 ( .gnd(gnd), .vdd(vdd), .A(_10697_), .B(bloque_datos_48_bF_buf1_), .Y(_10719_) );
NAND2X1 NAND2X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_10708_), .B(_10719_), .Y(_10730_) );
NAND2X1 NAND2X1_1550 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_64_bF_buf2_), .B(_10730_), .Y(_10741_) );
OR2X2 OR2X2_263 ( .gnd(gnd), .vdd(vdd), .A(_10730_), .B(bloque_datos_64_bF_buf1_), .Y(_10752_) );
NAND2X1 NAND2X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_10741_), .B(_10752_), .Y(_10763_) );
NAND2X1 NAND2X1_1552 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf1_), .B(_10763_), .Y(_10774_) );
OR2X2 OR2X2_264 ( .gnd(gnd), .vdd(vdd), .A(_10763_), .B(bloque_datos_80_bF_buf0_), .Y(_10785_) );
NAND2X1 NAND2X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_10774_), .B(_10785_), .Y(_10796_) );
NAND2X1 NAND2X1_1554 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_128_), .B(_10796_), .Y(_10807_) );
OR2X2 OR2X2_265 ( .gnd(gnd), .vdd(vdd), .A(_10796_), .B(module_2_W_128_), .Y(_10818_) );
NAND2X1 NAND2X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_10807_), .B(_10818_), .Y(_10829_) );
NAND2X1 NAND2X1_1556 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_144_), .B(_10829_), .Y(_10840_) );
OR2X2 OR2X2_266 ( .gnd(gnd), .vdd(vdd), .A(_10829_), .B(module_2_W_144_), .Y(_10851_) );
NAND2X1 NAND2X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_10840_), .B(_10851_), .Y(_10862_) );
NAND2X1 NAND2X1_1558 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_160_), .B(_10862_), .Y(_10873_) );
OR2X2 OR2X2_267 ( .gnd(gnd), .vdd(vdd), .A(_10862_), .B(module_2_W_160_), .Y(_10884_) );
NAND2X1 NAND2X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_10873_), .B(_10884_), .Y(_10895_) );
NAND2X1 NAND2X1_1560 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_176_), .B(_10895_), .Y(_10906_) );
OR2X2 OR2X2_268 ( .gnd(gnd), .vdd(vdd), .A(_10895_), .B(module_2_W_176_), .Y(_10917_) );
NAND2X1 NAND2X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_10906_), .B(_10917_), .Y(_10928_) );
NAND2X1 NAND2X1_1562 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_192_), .B(_10928_), .Y(_10939_) );
OR2X2 OR2X2_269 ( .gnd(gnd), .vdd(vdd), .A(_10928_), .B(module_2_W_192_), .Y(_10950_) );
NAND2X1 NAND2X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_10939_), .B(_10950_), .Y(_10961_) );
NAND2X1 NAND2X1_1564 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_208_), .B(_10961_), .Y(_10972_) );
OR2X2 OR2X2_270 ( .gnd(gnd), .vdd(vdd), .A(_10961_), .B(module_2_W_208_), .Y(_10983_) );
NAND2X1 NAND2X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_10972_), .B(_10983_), .Y(_10994_) );
INVX2 INVX2_382 ( .gnd(gnd), .vdd(vdd), .A(_10994_), .Y(_11005_) );
NOR2X1 NOR2X1_877 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_224_), .B(_11005_), .Y(_11016_) );
INVX1 INVX1_1625 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_225_), .Y(_11027_) );
INVX2 INVX2_383 ( .gnd(gnd), .vdd(vdd), .A(_10961_), .Y(_11038_) );
NOR2X1 NOR2X1_878 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_208_), .B(_11038_), .Y(_11049_) );
INVX2 INVX2_384 ( .gnd(gnd), .vdd(vdd), .A(_10928_), .Y(_11059_) );
NOR2X1 NOR2X1_879 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_192_), .B(_11059_), .Y(_11070_) );
INVX1 INVX1_1626 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_193_), .Y(_11081_) );
INVX2 INVX2_385 ( .gnd(gnd), .vdd(vdd), .A(_10895_), .Y(_11092_) );
NOR2X1 NOR2X1_880 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_176_), .B(_11092_), .Y(_11103_) );
INVX2 INVX2_386 ( .gnd(gnd), .vdd(vdd), .A(_10862_), .Y(_11114_) );
NOR2X1 NOR2X1_881 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_160_), .B(_11114_), .Y(_11125_) );
INVX1 INVX1_1627 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_161_), .Y(_11136_) );
INVX2 INVX2_387 ( .gnd(gnd), .vdd(vdd), .A(_10829_), .Y(_11147_) );
NOR2X1 NOR2X1_882 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_144_), .B(_11147_), .Y(_11158_) );
INVX1 INVX1_1628 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_145_), .Y(_11169_) );
INVX2 INVX2_388 ( .gnd(gnd), .vdd(vdd), .A(_10796_), .Y(_11180_) );
NOR2X1 NOR2X1_883 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_128_), .B(_11180_), .Y(_11191_) );
INVX2 INVX2_389 ( .gnd(gnd), .vdd(vdd), .A(_10763_), .Y(_11202_) );
NOR2X1 NOR2X1_884 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf5_), .B(_11202_), .Y(_11213_) );
AOI21X1 AOI21X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_10708_), .B(_10719_), .C(bloque_datos_64_bF_buf0_), .Y(_11224_) );
AOI21X1 AOI21X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_10676_), .B(_10686_), .C(bloque_datos_48_bF_buf0_), .Y(_11235_) );
INVX1 INVX1_1629 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_49_bF_buf3_), .Y(_11246_) );
AOI21X1 AOI21X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_10647_), .B(_10658_), .C(bloque_datos_32_bF_buf0_), .Y(_11257_) );
INVX1 INVX1_1630 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf1_), .Y(_11268_) );
AOI21X1 AOI21X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_10592_), .B(_10625_), .C(bloque_datos_16_bF_buf1_), .Y(_11279_) );
OAI21X1 OAI21X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_10570_), .B(_10581_), .C(_10603_), .Y(_11290_) );
INVX1 INVX1_1631 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(_11301_) );
INVX2 INVX2_390 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_0_), .Y(_11312_) );
NOR2X1 NOR2X1_885 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_16_), .B(_11312_), .Y(_11323_) );
NAND2X1 NAND2X1_1566 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_0_), .B(module_2_W_1_), .Y(_11334_) );
OR2X2 OR2X2_271 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_0_), .B(module_2_W_1_), .Y(_11345_) );
AOI21X1 AOI21X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_11334_), .B(_11345_), .C(module_2_W_17_), .Y(_11356_) );
INVX1 INVX1_1632 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_17_), .Y(_11367_) );
AND2X2 AND2X2_257 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_0_), .B(module_2_W_1_), .Y(_11378_) );
NOR2X1 NOR2X1_886 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_0_), .B(module_2_W_1_), .Y(_11389_) );
NOR3X1 NOR3X1_338 ( .gnd(gnd), .vdd(vdd), .A(_11367_), .B(_11389_), .C(_11378_), .Y(_11400_) );
OAI21X1 OAI21X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_11400_), .B(_11356_), .C(_11323_), .Y(_11411_) );
INVX1 INVX1_1633 ( .gnd(gnd), .vdd(vdd), .A(_11323_), .Y(_11421_) );
OAI21X1 OAI21X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_11378_), .B(_11389_), .C(_11367_), .Y(_11432_) );
NAND3X1 NAND3X1_2762 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_17_), .B(_11334_), .C(_11345_), .Y(_11443_) );
NAND3X1 NAND3X1_2763 ( .gnd(gnd), .vdd(vdd), .A(_11432_), .B(_11443_), .C(_11421_), .Y(_11454_) );
NAND2X1 NAND2X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_11454_), .B(_11411_), .Y(_11465_) );
NAND2X1 NAND2X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_11301_), .B(_11465_), .Y(_11476_) );
OR2X2 OR2X2_272 ( .gnd(gnd), .vdd(vdd), .A(_11465_), .B(_11301_), .Y(_11487_) );
NAND2X1 NAND2X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_11476_), .B(_11487_), .Y(_11498_) );
XNOR2X1 XNOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_11498_), .B(_11290_), .Y(_11509_) );
XNOR2X1 XNOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_11509_), .B(bloque_datos[17]), .Y(_11520_) );
AND2X2 AND2X2_258 ( .gnd(gnd), .vdd(vdd), .A(_11520_), .B(_11279_), .Y(_11531_) );
NOR2X1 NOR2X1_887 ( .gnd(gnd), .vdd(vdd), .A(_11279_), .B(_11520_), .Y(_11542_) );
OAI21X1 OAI21X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_11531_), .B(_11542_), .C(_11268_), .Y(_11553_) );
OR2X2 OR2X2_273 ( .gnd(gnd), .vdd(vdd), .A(_11531_), .B(_11542_), .Y(_11564_) );
NOR2X1 NOR2X1_888 ( .gnd(gnd), .vdd(vdd), .A(_11268_), .B(_11564_), .Y(_11575_) );
INVX1 INVX1_1634 ( .gnd(gnd), .vdd(vdd), .A(_11575_), .Y(_11586_) );
NAND2X1 NAND2X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_11553_), .B(_11586_), .Y(_11597_) );
AND2X2 AND2X2_259 ( .gnd(gnd), .vdd(vdd), .A(_11597_), .B(_11257_), .Y(_11608_) );
NOR2X1 NOR2X1_889 ( .gnd(gnd), .vdd(vdd), .A(_11257_), .B(_11597_), .Y(_11619_) );
OAI21X1 OAI21X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_11608_), .B(_11619_), .C(_11246_), .Y(_11630_) );
OR2X2 OR2X2_274 ( .gnd(gnd), .vdd(vdd), .A(_11608_), .B(_11619_), .Y(_11641_) );
NOR2X1 NOR2X1_890 ( .gnd(gnd), .vdd(vdd), .A(_11246_), .B(_11641_), .Y(_11652_) );
INVX1 INVX1_1635 ( .gnd(gnd), .vdd(vdd), .A(_11652_), .Y(_11663_) );
NAND2X1 NAND2X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_11630_), .B(_11663_), .Y(_11674_) );
AND2X2 AND2X2_260 ( .gnd(gnd), .vdd(vdd), .A(_11674_), .B(_11235_), .Y(_11685_) );
NOR2X1 NOR2X1_891 ( .gnd(gnd), .vdd(vdd), .A(_11235_), .B(_11674_), .Y(_11696_) );
NOR2X1 NOR2X1_892 ( .gnd(gnd), .vdd(vdd), .A(_11696_), .B(_11685_), .Y(_11707_) );
XNOR2X1 XNOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_11707_), .B(bloque_datos_65_bF_buf1_), .Y(_11718_) );
AND2X2 AND2X2_261 ( .gnd(gnd), .vdd(vdd), .A(_11718_), .B(_11224_), .Y(_11729_) );
NOR2X1 NOR2X1_893 ( .gnd(gnd), .vdd(vdd), .A(_11224_), .B(_11718_), .Y(_11740_) );
NOR2X1 NOR2X1_894 ( .gnd(gnd), .vdd(vdd), .A(_11740_), .B(_11729_), .Y(_11751_) );
NOR2X1 NOR2X1_895 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf2_), .B(_11751_), .Y(_11761_) );
INVX1 INVX1_1636 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf1_), .Y(_11772_) );
INVX1 INVX1_1637 ( .gnd(gnd), .vdd(vdd), .A(_11751_), .Y(_11783_) );
NOR2X1 NOR2X1_896 ( .gnd(gnd), .vdd(vdd), .A(_11772_), .B(_11783_), .Y(_11794_) );
OAI21X1 OAI21X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_11794_), .B(_11761_), .C(_11213_), .Y(_11805_) );
OR2X2 OR2X2_275 ( .gnd(gnd), .vdd(vdd), .A(_11794_), .B(_11761_), .Y(_11816_) );
NOR2X1 NOR2X1_897 ( .gnd(gnd), .vdd(vdd), .A(_11213_), .B(_11816_), .Y(_11827_) );
INVX2 INVX2_391 ( .gnd(gnd), .vdd(vdd), .A(_11827_), .Y(_11838_) );
NAND2X1 NAND2X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_11805_), .B(_11838_), .Y(_11849_) );
INVX2 INVX2_392 ( .gnd(gnd), .vdd(vdd), .A(_11849_), .Y(_11860_) );
NOR2X1 NOR2X1_898 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_129_), .B(_11860_), .Y(_11871_) );
AND2X2 AND2X2_262 ( .gnd(gnd), .vdd(vdd), .A(_11860_), .B(module_2_W_129_), .Y(_11882_) );
OAI21X1 OAI21X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_11882_), .B(_11871_), .C(_11191_), .Y(_11893_) );
OR2X2 OR2X2_276 ( .gnd(gnd), .vdd(vdd), .A(_11882_), .B(_11871_), .Y(_11904_) );
OR2X2 OR2X2_277 ( .gnd(gnd), .vdd(vdd), .A(_11904_), .B(_11191_), .Y(_11915_) );
NAND2X1 NAND2X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_11893_), .B(_11915_), .Y(_11926_) );
NAND2X1 NAND2X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_11169_), .B(_11926_), .Y(_11937_) );
NOR2X1 NOR2X1_899 ( .gnd(gnd), .vdd(vdd), .A(_11169_), .B(_11926_), .Y(_11948_) );
INVX1 INVX1_1638 ( .gnd(gnd), .vdd(vdd), .A(_11948_), .Y(_11959_) );
NAND2X1 NAND2X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_11937_), .B(_11959_), .Y(_11970_) );
NAND2X1 NAND2X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .B(_11970_), .Y(_11981_) );
NOR2X1 NOR2X1_900 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .B(_11970_), .Y(_11992_) );
INVX1 INVX1_1639 ( .gnd(gnd), .vdd(vdd), .A(_11992_), .Y(_12003_) );
NAND2X1 NAND2X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_11981_), .B(_12003_), .Y(_12010_) );
NAND2X1 NAND2X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_11136_), .B(_12010_), .Y(_12011_) );
NOR2X1 NOR2X1_901 ( .gnd(gnd), .vdd(vdd), .A(_11136_), .B(_12010_), .Y(_12012_) );
INVX1 INVX1_1640 ( .gnd(gnd), .vdd(vdd), .A(_12012_), .Y(_12013_) );
NAND2X1 NAND2X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_12011_), .B(_12013_), .Y(_12014_) );
NAND2X1 NAND2X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_11125_), .B(_12014_), .Y(_12015_) );
NOR2X1 NOR2X1_902 ( .gnd(gnd), .vdd(vdd), .A(_11125_), .B(_12014_), .Y(_12016_) );
INVX1 INVX1_1641 ( .gnd(gnd), .vdd(vdd), .A(_12016_), .Y(_12017_) );
NAND2X1 NAND2X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_12015_), .B(_12017_), .Y(_12018_) );
INVX2 INVX2_393 ( .gnd(gnd), .vdd(vdd), .A(_12018_), .Y(_12019_) );
NOR2X1 NOR2X1_903 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_177_), .B(_12019_), .Y(_12020_) );
NAND2X1 NAND2X1_1582 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_177_), .B(_12019_), .Y(_12021_) );
INVX2 INVX2_394 ( .gnd(gnd), .vdd(vdd), .A(_12021_), .Y(_12022_) );
OAI21X1 OAI21X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_12022_), .B(_12020_), .C(_11103_), .Y(_12023_) );
OR2X2 OR2X2_278 ( .gnd(gnd), .vdd(vdd), .A(_12022_), .B(_12020_), .Y(_12024_) );
NOR2X1 NOR2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_11103_), .B(_12024_), .Y(_12025_) );
INVX1 INVX1_1642 ( .gnd(gnd), .vdd(vdd), .A(_12025_), .Y(_12026_) );
NAND2X1 NAND2X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_12023_), .B(_12026_), .Y(_12027_) );
NAND2X1 NAND2X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_11081_), .B(_12027_), .Y(_12028_) );
NOR2X1 NOR2X1_905 ( .gnd(gnd), .vdd(vdd), .A(_11081_), .B(_12027_), .Y(_12029_) );
INVX1 INVX1_1643 ( .gnd(gnd), .vdd(vdd), .A(_12029_), .Y(_12030_) );
NAND2X1 NAND2X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_12028_), .B(_12030_), .Y(_12031_) );
NAND2X1 NAND2X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_11070_), .B(_12031_), .Y(_12032_) );
NOR2X1 NOR2X1_906 ( .gnd(gnd), .vdd(vdd), .A(_11070_), .B(_12031_), .Y(_12033_) );
INVX1 INVX1_1644 ( .gnd(gnd), .vdd(vdd), .A(_12033_), .Y(_12034_) );
NAND2X1 NAND2X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_12032_), .B(_12034_), .Y(_12035_) );
INVX2 INVX2_395 ( .gnd(gnd), .vdd(vdd), .A(_12035_), .Y(_12036_) );
NOR2X1 NOR2X1_907 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_209_), .B(_12036_), .Y(_12037_) );
NAND2X1 NAND2X1_1588 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_209_), .B(_12036_), .Y(_12038_) );
INVX2 INVX2_396 ( .gnd(gnd), .vdd(vdd), .A(_12038_), .Y(_12039_) );
OAI21X1 OAI21X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_12039_), .B(_12037_), .C(_11049_), .Y(_12040_) );
OR2X2 OR2X2_279 ( .gnd(gnd), .vdd(vdd), .A(_12039_), .B(_12037_), .Y(_12041_) );
NOR2X1 NOR2X1_908 ( .gnd(gnd), .vdd(vdd), .A(_11049_), .B(_12041_), .Y(_12042_) );
INVX2 INVX2_397 ( .gnd(gnd), .vdd(vdd), .A(_12042_), .Y(_12043_) );
NAND2X1 NAND2X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_12040_), .B(_12043_), .Y(_12044_) );
NAND2X1 NAND2X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_11027_), .B(_12044_), .Y(_12045_) );
NOR2X1 NOR2X1_909 ( .gnd(gnd), .vdd(vdd), .A(_11027_), .B(_12044_), .Y(_12046_) );
INVX1 INVX1_1645 ( .gnd(gnd), .vdd(vdd), .A(_12046_), .Y(_12047_) );
NAND2X1 NAND2X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_12045_), .B(_12047_), .Y(_12048_) );
NAND2X1 NAND2X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_11016_), .B(_12048_), .Y(_12049_) );
NOR2X1 NOR2X1_910 ( .gnd(gnd), .vdd(vdd), .A(_11016_), .B(_12048_), .Y(_12050_) );
INVX1 INVX1_1646 ( .gnd(gnd), .vdd(vdd), .A(_12050_), .Y(_12051_) );
NAND2X1 NAND2X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_12049_), .B(_12051_), .Y(_12052_) );
NOR2X1 NOR2X1_911 ( .gnd(gnd), .vdd(vdd), .A(_10559_), .B(_12052_), .Y(_12053_) );
INVX1 INVX1_1647 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_242_), .Y(_12054_) );
INVX1 INVX1_1648 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_194_), .Y(_12055_) );
INVX1 INVX1_1649 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_178_), .Y(_12056_) );
INVX1 INVX1_1650 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_162_), .Y(_12057_) );
NOR2X1 NOR2X1_912 ( .gnd(gnd), .vdd(vdd), .A(_11191_), .B(_11904_), .Y(_12058_) );
AND2X2 AND2X2_263 ( .gnd(gnd), .vdd(vdd), .A(_11707_), .B(bloque_datos_65_bF_buf0_), .Y(_12059_) );
INVX1 INVX1_1651 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf2_), .Y(_12060_) );
INVX1 INVX1_1652 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf2_), .Y(_12061_) );
INVX1 INVX1_1653 ( .gnd(gnd), .vdd(vdd), .A(_11542_), .Y(_12062_) );
NAND2X1 NAND2X1_1594 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .B(_11509_), .Y(_12063_) );
INVX1 INVX1_1654 ( .gnd(gnd), .vdd(vdd), .A(_11290_), .Y(_12064_) );
NOR2X1 NOR2X1_913 ( .gnd(gnd), .vdd(vdd), .A(_12064_), .B(_11498_), .Y(_12065_) );
INVX1 INVX1_1655 ( .gnd(gnd), .vdd(vdd), .A(_11487_), .Y(_12066_) );
INVX1 INVX1_1656 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf3_), .Y(_12067_) );
INVX1 INVX1_1657 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_18_), .Y(_12068_) );
NAND3X1 NAND3X1_2764 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_2_), .B(module_2_W_0_), .C(module_2_W_1_), .Y(_12069_) );
INVX2 INVX2_398 ( .gnd(gnd), .vdd(vdd), .A(_12069_), .Y(_12070_) );
AOI21X1 AOI21X1_1674 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_0_), .B(module_2_W_1_), .C(module_2_W_2_), .Y(_12071_) );
OAI21X1 OAI21X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_12070_), .B(_12071_), .C(_12068_), .Y(_12072_) );
INVX2 INVX2_399 ( .gnd(gnd), .vdd(vdd), .A(_12071_), .Y(_12073_) );
NAND3X1 NAND3X1_2765 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_18_), .B(_12069_), .C(_12073_), .Y(_12074_) );
NAND3X1 NAND3X1_2766 ( .gnd(gnd), .vdd(vdd), .A(_11400_), .B(_12074_), .C(_12072_), .Y(_12075_) );
AOI21X1 AOI21X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_12069_), .B(_12073_), .C(module_2_W_18_), .Y(_12076_) );
NOR3X1 NOR3X1_339 ( .gnd(gnd), .vdd(vdd), .A(_12068_), .B(_12071_), .C(_12070_), .Y(_12077_) );
OAI21X1 OAI21X1_1904 ( .gnd(gnd), .vdd(vdd), .A(_12077_), .B(_12076_), .C(_11443_), .Y(_12078_) );
NAND2X1 NAND2X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_12075_), .B(_12078_), .Y(_12079_) );
NOR2X1 NOR2X1_914 ( .gnd(gnd), .vdd(vdd), .A(_11454_), .B(_12079_), .Y(_12080_) );
INVX1 INVX1_1658 ( .gnd(gnd), .vdd(vdd), .A(_11454_), .Y(_12081_) );
AOI21X1 AOI21X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_12075_), .B(_12078_), .C(_12081_), .Y(_12082_) );
OAI21X1 OAI21X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_12080_), .B(_12082_), .C(_12067_), .Y(_12083_) );
OR2X2 OR2X2_280 ( .gnd(gnd), .vdd(vdd), .A(_12079_), .B(_11454_), .Y(_12084_) );
INVX1 INVX1_1659 ( .gnd(gnd), .vdd(vdd), .A(_12082_), .Y(_12085_) );
NAND3X1 NAND3X1_2767 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf2_), .B(_12085_), .C(_12084_), .Y(_12086_) );
NAND3X1 NAND3X1_2768 ( .gnd(gnd), .vdd(vdd), .A(_12066_), .B(_12083_), .C(_12086_), .Y(_12087_) );
AOI21X1 AOI21X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_12085_), .B(_12084_), .C(bloque_datos_2_bF_buf1_), .Y(_12088_) );
NOR3X1 NOR3X1_340 ( .gnd(gnd), .vdd(vdd), .A(_12067_), .B(_12082_), .C(_12080_), .Y(_12089_) );
OAI21X1 OAI21X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_12088_), .B(_12089_), .C(_11487_), .Y(_12090_) );
NAND3X1 NAND3X1_2769 ( .gnd(gnd), .vdd(vdd), .A(_12065_), .B(_12087_), .C(_12090_), .Y(_12091_) );
AOI21X1 AOI21X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_12087_), .B(_12090_), .C(_12065_), .Y(_12092_) );
INVX1 INVX1_1660 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .Y(_12093_) );
AOI21X1 AOI21X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_12091_), .B(_12093_), .C(bloque_datos[18]), .Y(_12094_) );
INVX1 INVX1_1661 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .Y(_12095_) );
INVX1 INVX1_1662 ( .gnd(gnd), .vdd(vdd), .A(_12065_), .Y(_12096_) );
NOR3X1 NOR3X1_341 ( .gnd(gnd), .vdd(vdd), .A(_12089_), .B(_11487_), .C(_12088_), .Y(_12097_) );
AOI21X1 AOI21X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_12083_), .B(_12086_), .C(_12066_), .Y(_12098_) );
NOR3X1 NOR3X1_342 ( .gnd(gnd), .vdd(vdd), .A(_12096_), .B(_12098_), .C(_12097_), .Y(_12099_) );
NOR3X1 NOR3X1_343 ( .gnd(gnd), .vdd(vdd), .A(_12095_), .B(_12092_), .C(_12099_), .Y(_12100_) );
NOR3X1 NOR3X1_344 ( .gnd(gnd), .vdd(vdd), .A(_12063_), .B(_12100_), .C(_12094_), .Y(_12101_) );
INVX1 INVX1_1663 ( .gnd(gnd), .vdd(vdd), .A(_12063_), .Y(_12102_) );
OAI21X1 OAI21X1_1907 ( .gnd(gnd), .vdd(vdd), .A(_12099_), .B(_12092_), .C(_12095_), .Y(_12103_) );
INVX2 INVX2_400 ( .gnd(gnd), .vdd(vdd), .A(_12100_), .Y(_12104_) );
AOI21X1 AOI21X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_12103_), .B(_12104_), .C(_12102_), .Y(_12105_) );
NOR3X1 NOR3X1_345 ( .gnd(gnd), .vdd(vdd), .A(_12062_), .B(_12101_), .C(_12105_), .Y(_12106_) );
NAND3X1 NAND3X1_2770 ( .gnd(gnd), .vdd(vdd), .A(_12102_), .B(_12103_), .C(_12104_), .Y(_12107_) );
OAI21X1 OAI21X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_12094_), .B(_12100_), .C(_12063_), .Y(_12108_) );
AOI21X1 AOI21X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_12108_), .B(_12107_), .C(_11542_), .Y(_12109_) );
OAI21X1 OAI21X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_12106_), .B(_12109_), .C(_12061_), .Y(_12110_) );
NAND3X1 NAND3X1_2771 ( .gnd(gnd), .vdd(vdd), .A(_11542_), .B(_12108_), .C(_12107_), .Y(_12111_) );
OAI21X1 OAI21X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_12105_), .B(_12101_), .C(_12062_), .Y(_12112_) );
NAND3X1 NAND3X1_2772 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf1_), .B(_12111_), .C(_12112_), .Y(_12113_) );
NAND3X1 NAND3X1_2773 ( .gnd(gnd), .vdd(vdd), .A(_11575_), .B(_12113_), .C(_12110_), .Y(_12114_) );
AOI21X1 AOI21X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_12111_), .B(_12112_), .C(bloque_datos_34_bF_buf0_), .Y(_12115_) );
NOR3X1 NOR3X1_346 ( .gnd(gnd), .vdd(vdd), .A(_12061_), .B(_12109_), .C(_12106_), .Y(_12116_) );
OAI21X1 OAI21X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_12116_), .B(_12115_), .C(_11586_), .Y(_12117_) );
NAND3X1 NAND3X1_2774 ( .gnd(gnd), .vdd(vdd), .A(_11619_), .B(_12114_), .C(_12117_), .Y(_12118_) );
AOI21X1 AOI21X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_12114_), .B(_12117_), .C(_11619_), .Y(_12119_) );
INVX1 INVX1_1664 ( .gnd(gnd), .vdd(vdd), .A(_12119_), .Y(_12120_) );
AOI21X1 AOI21X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_12118_), .B(_12120_), .C(bloque_datos_50_bF_buf1_), .Y(_12121_) );
INVX1 INVX1_1665 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_50_bF_buf0_), .Y(_12122_) );
INVX1 INVX1_1666 ( .gnd(gnd), .vdd(vdd), .A(_12118_), .Y(_12123_) );
NOR3X1 NOR3X1_347 ( .gnd(gnd), .vdd(vdd), .A(_12122_), .B(_12119_), .C(_12123_), .Y(_12124_) );
NOR2X1 NOR2X1_915 ( .gnd(gnd), .vdd(vdd), .A(_12121_), .B(_12124_), .Y(_12125_) );
NAND2X1 NAND2X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_11652_), .B(_12125_), .Y(_12126_) );
OAI21X1 OAI21X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_12124_), .B(_12121_), .C(_11663_), .Y(_12127_) );
NAND3X1 NAND3X1_2775 ( .gnd(gnd), .vdd(vdd), .A(_11696_), .B(_12127_), .C(_12126_), .Y(_12128_) );
INVX2 INVX2_401 ( .gnd(gnd), .vdd(vdd), .A(_12128_), .Y(_12129_) );
AOI21X1 AOI21X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_12127_), .B(_12126_), .C(_11696_), .Y(_12130_) );
OAI21X1 OAI21X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_12129_), .B(_12130_), .C(_12060_), .Y(_12131_) );
INVX1 INVX1_1667 ( .gnd(gnd), .vdd(vdd), .A(_11696_), .Y(_12132_) );
AND2X2 AND2X2_264 ( .gnd(gnd), .vdd(vdd), .A(_12125_), .B(_11652_), .Y(_12133_) );
INVX1 INVX1_1668 ( .gnd(gnd), .vdd(vdd), .A(_12127_), .Y(_12134_) );
OAI21X1 OAI21X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_12133_), .B(_12134_), .C(_12132_), .Y(_12135_) );
NAND3X1 NAND3X1_2776 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf1_), .B(_12128_), .C(_12135_), .Y(_12136_) );
NAND3X1 NAND3X1_2777 ( .gnd(gnd), .vdd(vdd), .A(_12059_), .B(_12136_), .C(_12131_), .Y(_12137_) );
INVX1 INVX1_1669 ( .gnd(gnd), .vdd(vdd), .A(_12059_), .Y(_12138_) );
AOI21X1 AOI21X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_12128_), .B(_12135_), .C(bloque_datos_66_bF_buf0_), .Y(_12139_) );
NOR3X1 NOR3X1_348 ( .gnd(gnd), .vdd(vdd), .A(_12060_), .B(_12130_), .C(_12129_), .Y(_12140_) );
OAI21X1 OAI21X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_12140_), .B(_12139_), .C(_12138_), .Y(_12141_) );
NAND3X1 NAND3X1_2778 ( .gnd(gnd), .vdd(vdd), .A(_11740_), .B(_12137_), .C(_12141_), .Y(_12142_) );
INVX2 INVX2_402 ( .gnd(gnd), .vdd(vdd), .A(_11740_), .Y(_12143_) );
NOR3X1 NOR3X1_349 ( .gnd(gnd), .vdd(vdd), .A(_12138_), .B(_12139_), .C(_12140_), .Y(_12144_) );
AOI21X1 AOI21X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_12136_), .B(_12131_), .C(_12059_), .Y(_12145_) );
OAI21X1 OAI21X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_12144_), .B(_12145_), .C(_12143_), .Y(_12146_) );
AOI21X1 AOI21X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_12142_), .B(_12146_), .C(bloque_datos_82_bF_buf0_), .Y(_12147_) );
INVX1 INVX1_1670 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf4_), .Y(_12148_) );
NOR3X1 NOR3X1_350 ( .gnd(gnd), .vdd(vdd), .A(_12143_), .B(_12145_), .C(_12144_), .Y(_12149_) );
AOI21X1 AOI21X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_12137_), .B(_12141_), .C(_11740_), .Y(_12150_) );
NOR3X1 NOR3X1_351 ( .gnd(gnd), .vdd(vdd), .A(_12148_), .B(_12150_), .C(_12149_), .Y(_12151_) );
NOR2X1 NOR2X1_916 ( .gnd(gnd), .vdd(vdd), .A(_12147_), .B(_12151_), .Y(_12152_) );
NAND2X1 NAND2X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_11794_), .B(_12152_), .Y(_12153_) );
OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_11772_), .B(_11783_), .C(_12151_), .D(_12147_), .Y(_12154_) );
NAND3X1 NAND3X1_2779 ( .gnd(gnd), .vdd(vdd), .A(_11827_), .B(_12154_), .C(_12153_), .Y(_12155_) );
AND2X2 AND2X2_265 ( .gnd(gnd), .vdd(vdd), .A(_12152_), .B(_11794_), .Y(_12156_) );
INVX2 INVX2_403 ( .gnd(gnd), .vdd(vdd), .A(_12154_), .Y(_12157_) );
OAI21X1 OAI21X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_12156_), .B(_12157_), .C(_11838_), .Y(_12158_) );
AOI21X1 AOI21X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_12155_), .B(_12158_), .C(module_2_W_130_), .Y(_12159_) );
INVX1 INVX1_1671 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_130_), .Y(_12160_) );
NOR3X1 NOR3X1_352 ( .gnd(gnd), .vdd(vdd), .A(_12157_), .B(_11838_), .C(_12156_), .Y(_12161_) );
AOI21X1 AOI21X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_12154_), .B(_12153_), .C(_11827_), .Y(_12162_) );
NOR3X1 NOR3X1_353 ( .gnd(gnd), .vdd(vdd), .A(_12160_), .B(_12162_), .C(_12161_), .Y(_12163_) );
NOR2X1 NOR2X1_917 ( .gnd(gnd), .vdd(vdd), .A(_12159_), .B(_12163_), .Y(_12164_) );
NAND2X1 NAND2X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_11882_), .B(_12164_), .Y(_12165_) );
NOR2X1 NOR2X1_918 ( .gnd(gnd), .vdd(vdd), .A(_11882_), .B(_12164_), .Y(_12166_) );
INVX1 INVX1_1672 ( .gnd(gnd), .vdd(vdd), .A(_12166_), .Y(_12167_) );
NAND3X1 NAND3X1_2780 ( .gnd(gnd), .vdd(vdd), .A(_12058_), .B(_12165_), .C(_12167_), .Y(_12168_) );
INVX1 INVX1_1673 ( .gnd(gnd), .vdd(vdd), .A(_12165_), .Y(_12169_) );
OAI21X1 OAI21X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_12169_), .B(_12166_), .C(_11915_), .Y(_12170_) );
AOI21X1 AOI21X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_12170_), .B(_12168_), .C(module_2_W_146_), .Y(_12171_) );
INVX1 INVX1_1674 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_146_), .Y(_12172_) );
NOR3X1 NOR3X1_354 ( .gnd(gnd), .vdd(vdd), .A(_11915_), .B(_12166_), .C(_12169_), .Y(_12173_) );
AOI21X1 AOI21X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_12165_), .B(_12167_), .C(_12058_), .Y(_12174_) );
NOR3X1 NOR3X1_355 ( .gnd(gnd), .vdd(vdd), .A(_12173_), .B(_12172_), .C(_12174_), .Y(_12175_) );
NOR2X1 NOR2X1_919 ( .gnd(gnd), .vdd(vdd), .A(_12171_), .B(_12175_), .Y(_12176_) );
NAND2X1 NAND2X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_11948_), .B(_12176_), .Y(_12177_) );
OAI21X1 OAI21X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_12175_), .B(_12171_), .C(_11959_), .Y(_12178_) );
AND2X2 AND2X2_266 ( .gnd(gnd), .vdd(vdd), .A(_12177_), .B(_12178_), .Y(_12179_) );
NAND2X1 NAND2X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_11992_), .B(_12179_), .Y(_12180_) );
INVX1 INVX1_1675 ( .gnd(gnd), .vdd(vdd), .A(_12180_), .Y(_12181_) );
NOR2X1 NOR2X1_920 ( .gnd(gnd), .vdd(vdd), .A(_11992_), .B(_12179_), .Y(_12182_) );
OAI21X1 OAI21X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_12181_), .B(_12182_), .C(_12057_), .Y(_12183_) );
NOR2X1 NOR2X1_921 ( .gnd(gnd), .vdd(vdd), .A(_12182_), .B(_12181_), .Y(_12184_) );
NAND2X1 NAND2X1_1601 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_162_), .B(_12184_), .Y(_12185_) );
NAND3X1 NAND3X1_2781 ( .gnd(gnd), .vdd(vdd), .A(_12012_), .B(_12183_), .C(_12185_), .Y(_12186_) );
INVX1 INVX1_1676 ( .gnd(gnd), .vdd(vdd), .A(_12183_), .Y(_12187_) );
AND2X2 AND2X2_267 ( .gnd(gnd), .vdd(vdd), .A(_12184_), .B(module_2_W_162_), .Y(_12188_) );
OAI21X1 OAI21X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_12188_), .B(_12187_), .C(_12013_), .Y(_12189_) );
NAND3X1 NAND3X1_2782 ( .gnd(gnd), .vdd(vdd), .A(_12016_), .B(_12186_), .C(_12189_), .Y(_12190_) );
INVX2 INVX2_404 ( .gnd(gnd), .vdd(vdd), .A(_12190_), .Y(_12191_) );
AOI21X1 AOI21X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_12186_), .B(_12189_), .C(_12016_), .Y(_12192_) );
OAI21X1 OAI21X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_12191_), .B(_12192_), .C(_12056_), .Y(_12193_) );
NOR2X1 NOR2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_12192_), .B(_12191_), .Y(_12194_) );
NAND2X1 NAND2X1_1602 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_178_), .B(_12194_), .Y(_12195_) );
NAND3X1 NAND3X1_2783 ( .gnd(gnd), .vdd(vdd), .A(_12022_), .B(_12193_), .C(_12195_), .Y(_12196_) );
INVX1 INVX1_1677 ( .gnd(gnd), .vdd(vdd), .A(_12193_), .Y(_12197_) );
INVX1 INVX1_1678 ( .gnd(gnd), .vdd(vdd), .A(_12195_), .Y(_12198_) );
OAI21X1 OAI21X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_12198_), .B(_12197_), .C(_12021_), .Y(_12199_) );
NAND3X1 NAND3X1_2784 ( .gnd(gnd), .vdd(vdd), .A(_12025_), .B(_12196_), .C(_12199_), .Y(_12200_) );
INVX2 INVX2_405 ( .gnd(gnd), .vdd(vdd), .A(_12200_), .Y(_12201_) );
AOI21X1 AOI21X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_12196_), .B(_12199_), .C(_12025_), .Y(_12202_) );
OAI21X1 OAI21X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_12201_), .B(_12202_), .C(_12055_), .Y(_12203_) );
INVX1 INVX1_1679 ( .gnd(gnd), .vdd(vdd), .A(_12203_), .Y(_12204_) );
NOR3X1 NOR3X1_356 ( .gnd(gnd), .vdd(vdd), .A(_12055_), .B(_12202_), .C(_12201_), .Y(_12205_) );
NOR2X1 NOR2X1_923 ( .gnd(gnd), .vdd(vdd), .A(_12205_), .B(_12204_), .Y(_12206_) );
NAND2X1 NAND2X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_12029_), .B(_12206_), .Y(_12207_) );
OAI21X1 OAI21X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_12204_), .B(_12205_), .C(_12030_), .Y(_12208_) );
NAND3X1 NAND3X1_2785 ( .gnd(gnd), .vdd(vdd), .A(_12033_), .B(_12208_), .C(_12207_), .Y(_12209_) );
INVX2 INVX2_406 ( .gnd(gnd), .vdd(vdd), .A(_12209_), .Y(_12210_) );
AOI21X1 AOI21X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_12208_), .B(_12207_), .C(_12033_), .Y(_12211_) );
NOR2X1 NOR2X1_924 ( .gnd(gnd), .vdd(vdd), .A(_12211_), .B(_12210_), .Y(_12212_) );
NOR2X1 NOR2X1_925 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_210_), .B(_12212_), .Y(_12213_) );
INVX1 INVX1_1680 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_210_), .Y(_12214_) );
NOR3X1 NOR3X1_357 ( .gnd(gnd), .vdd(vdd), .A(_12214_), .B(_12211_), .C(_12210_), .Y(_12215_) );
NOR2X1 NOR2X1_926 ( .gnd(gnd), .vdd(vdd), .A(_12215_), .B(_12213_), .Y(_12216_) );
NAND2X1 NAND2X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_12039_), .B(_12216_), .Y(_12217_) );
INVX1 INVX1_1681 ( .gnd(gnd), .vdd(vdd), .A(_12217_), .Y(_12218_) );
OAI21X1 OAI21X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_12213_), .B(_12215_), .C(_12038_), .Y(_12219_) );
INVX2 INVX2_407 ( .gnd(gnd), .vdd(vdd), .A(_12219_), .Y(_12220_) );
NOR2X1 NOR2X1_927 ( .gnd(gnd), .vdd(vdd), .A(_12220_), .B(_12218_), .Y(_12221_) );
NAND2X1 NAND2X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_12042_), .B(_12221_), .Y(_12222_) );
OAI21X1 OAI21X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_12218_), .B(_12220_), .C(_12043_), .Y(_12223_) );
AOI21X1 AOI21X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_12223_), .B(_12222_), .C(module_2_W_226_), .Y(_12224_) );
INVX1 INVX1_1682 ( .gnd(gnd), .vdd(vdd), .A(_12224_), .Y(_12225_) );
NAND3X1 NAND3X1_2786 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_226_), .B(_12223_), .C(_12222_), .Y(_12226_) );
NAND3X1 NAND3X1_2787 ( .gnd(gnd), .vdd(vdd), .A(_12046_), .B(_12226_), .C(_12225_), .Y(_12227_) );
INVX2 INVX2_408 ( .gnd(gnd), .vdd(vdd), .A(_12226_), .Y(_12228_) );
OAI21X1 OAI21X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_12228_), .B(_12224_), .C(_12047_), .Y(_12229_) );
NAND3X1 NAND3X1_2788 ( .gnd(gnd), .vdd(vdd), .A(_12050_), .B(_12229_), .C(_12227_), .Y(_12230_) );
INVX1 INVX1_1683 ( .gnd(gnd), .vdd(vdd), .A(_12230_), .Y(_12231_) );
AOI21X1 AOI21X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_12229_), .B(_12227_), .C(_12050_), .Y(_12232_) );
OAI21X1 OAI21X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_12231_), .B(_12232_), .C(_12054_), .Y(_12233_) );
NOR2X1 NOR2X1_928 ( .gnd(gnd), .vdd(vdd), .A(_12232_), .B(_12231_), .Y(_12234_) );
NAND2X1 NAND2X1_1606 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_242_), .B(_12234_), .Y(_12235_) );
NAND3X1 NAND3X1_2789 ( .gnd(gnd), .vdd(vdd), .A(_12053_), .B(_12233_), .C(_12235_), .Y(_12236_) );
NAND2X1 NAND2X1_1607 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_224_), .B(_10994_), .Y(_12237_) );
OR2X2 OR2X2_281 ( .gnd(gnd), .vdd(vdd), .A(_10994_), .B(module_2_W_224_), .Y(_12238_) );
NAND2X1 NAND2X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_12237_), .B(_12238_), .Y(_12239_) );
INVX4 INVX4_10 ( .gnd(gnd), .vdd(vdd), .A(_12239_), .Y(_12240_) );
INVX2 INVX2_409 ( .gnd(gnd), .vdd(vdd), .A(_12052_), .Y(_12241_) );
NOR2X1 NOR2X1_929 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_241_), .B(_12241_), .Y(_12242_) );
NOR2X1 NOR2X1_930 ( .gnd(gnd), .vdd(vdd), .A(_12053_), .B(_12242_), .Y(_12243_) );
OAI21X1 OAI21X1_1930 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_240_), .B(_12240_), .C(_12243_), .Y(_12244_) );
INVX1 INVX1_1684 ( .gnd(gnd), .vdd(vdd), .A(_12053_), .Y(_12245_) );
INVX1 INVX1_1685 ( .gnd(gnd), .vdd(vdd), .A(_12233_), .Y(_12246_) );
INVX1 INVX1_1686 ( .gnd(gnd), .vdd(vdd), .A(_12235_), .Y(_12247_) );
OAI21X1 OAI21X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_12247_), .B(_12246_), .C(_12245_), .Y(_12248_) );
INVX1 INVX1_1687 ( .gnd(gnd), .vdd(vdd), .A(_12248_), .Y(_12249_) );
OAI21X1 OAI21X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_12249_), .B(_12244_), .C(_12236_), .Y(_12250_) );
INVX1 INVX1_1688 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_243_), .Y(_12251_) );
NAND2X1 NAND2X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_12227_), .B(_12230_), .Y(_12252_) );
INVX1 INVX1_1689 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_227_), .Y(_12253_) );
OAI21X1 OAI21X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_12043_), .B(_12220_), .C(_12217_), .Y(_12254_) );
INVX1 INVX1_1690 ( .gnd(gnd), .vdd(vdd), .A(_12215_), .Y(_12255_) );
INVX1 INVX1_1691 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_211_), .Y(_12256_) );
INVX1 INVX1_1692 ( .gnd(gnd), .vdd(vdd), .A(_12207_), .Y(_12257_) );
AOI21X1 AOI21X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_12033_), .B(_12208_), .C(_12257_), .Y(_12258_) );
INVX1 INVX1_1693 ( .gnd(gnd), .vdd(vdd), .A(_12205_), .Y(_12259_) );
INVX1 INVX1_1694 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_195_), .Y(_12260_) );
AND2X2 AND2X2_268 ( .gnd(gnd), .vdd(vdd), .A(_12200_), .B(_12196_), .Y(_12261_) );
INVX1 INVX1_1695 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_179_), .Y(_12262_) );
INVX1 INVX1_1696 ( .gnd(gnd), .vdd(vdd), .A(_12186_), .Y(_12263_) );
INVX1 INVX1_1697 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_163_), .Y(_12264_) );
INVX1 INVX1_1698 ( .gnd(gnd), .vdd(vdd), .A(_12178_), .Y(_12265_) );
OAI21X1 OAI21X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_12003_), .B(_12265_), .C(_12177_), .Y(_12266_) );
INVX1 INVX1_1699 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_147_), .Y(_12267_) );
OAI21X1 OAI21X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_11915_), .B(_12166_), .C(_12165_), .Y(_12268_) );
INVX1 INVX1_1700 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_131_), .Y(_12269_) );
OAI21X1 OAI21X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_11838_), .B(_12157_), .C(_12153_), .Y(_12270_) );
OAI21X1 OAI21X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_12145_), .B(_12143_), .C(_12137_), .Y(_12271_) );
OAI21X1 OAI21X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_12134_), .B(_12132_), .C(_12126_), .Y(_12272_) );
INVX1 INVX1_1701 ( .gnd(gnd), .vdd(vdd), .A(_12124_), .Y(_12273_) );
AND2X2 AND2X2_269 ( .gnd(gnd), .vdd(vdd), .A(_12118_), .B(_12114_), .Y(_12274_) );
AOI21X1 AOI21X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_12108_), .B(_11542_), .C(_12101_), .Y(_12275_) );
INVX2 INVX2_410 ( .gnd(gnd), .vdd(vdd), .A(_12275_), .Y(_12276_) );
OAI21X1 OAI21X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_12098_), .B(_12096_), .C(_12087_), .Y(_12277_) );
NOR3X1 NOR3X1_358 ( .gnd(gnd), .vdd(vdd), .A(_12076_), .B(_11443_), .C(_12077_), .Y(_12278_) );
AOI21X1 AOI21X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_12081_), .B(_12078_), .C(_12278_), .Y(_12279_) );
INVX1 INVX1_1702 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_19_), .Y(_12280_) );
INVX2 INVX2_411 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_3_), .Y(_12281_) );
NOR2X1 NOR2X1_931 ( .gnd(gnd), .vdd(vdd), .A(_12281_), .B(_12069_), .Y(_12282_) );
AND2X2 AND2X2_270 ( .gnd(gnd), .vdd(vdd), .A(_12069_), .B(_12281_), .Y(_12283_) );
OAI21X1 OAI21X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_12283_), .B(_12282_), .C(_12280_), .Y(_12284_) );
NOR2X1 NOR2X1_932 ( .gnd(gnd), .vdd(vdd), .A(_12282_), .B(_12283_), .Y(_12285_) );
NAND2X1 NAND2X1_1610 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_19_), .B(_12285_), .Y(_12286_) );
AOI21X1 AOI21X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_12284_), .B(_12286_), .C(_12074_), .Y(_12287_) );
INVX1 INVX1_1703 ( .gnd(gnd), .vdd(vdd), .A(_12282_), .Y(_12288_) );
NAND2X1 NAND2X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_12281_), .B(_12069_), .Y(_12289_) );
AOI21X1 AOI21X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_12289_), .B(_12288_), .C(module_2_W_19_), .Y(_12290_) );
NOR3X1 NOR3X1_359 ( .gnd(gnd), .vdd(vdd), .A(_12282_), .B(_12280_), .C(_12283_), .Y(_12291_) );
NOR3X1 NOR3X1_360 ( .gnd(gnd), .vdd(vdd), .A(_12077_), .B(_12291_), .C(_12290_), .Y(_12292_) );
OAI21X1 OAI21X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_12287_), .B(_12292_), .C(_12279_), .Y(_12293_) );
NOR2X1 NOR2X1_933 ( .gnd(gnd), .vdd(vdd), .A(_12292_), .B(_12287_), .Y(_12294_) );
OAI21X1 OAI21X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_12080_), .B(_12278_), .C(_12294_), .Y(_12295_) );
AOI21X1 AOI21X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_12293_), .B(_12295_), .C(bloque_datos_3_bF_buf3_), .Y(_12296_) );
INVX1 INVX1_1704 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf2_), .Y(_12297_) );
INVX1 INVX1_1705 ( .gnd(gnd), .vdd(vdd), .A(_12293_), .Y(_12298_) );
AOI21X1 AOI21X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_12074_), .B(_12072_), .C(_11400_), .Y(_12299_) );
OAI21X1 OAI21X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_12299_), .B(_11454_), .C(_12075_), .Y(_12300_) );
AND2X2 AND2X2_271 ( .gnd(gnd), .vdd(vdd), .A(_12294_), .B(_12300_), .Y(_12301_) );
NOR3X1 NOR3X1_361 ( .gnd(gnd), .vdd(vdd), .A(_12298_), .B(_12297_), .C(_12301_), .Y(_12302_) );
OAI21X1 OAI21X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_12302_), .B(_12296_), .C(_12089_), .Y(_12303_) );
OAI21X1 OAI21X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_12301_), .B(_12298_), .C(_12297_), .Y(_12304_) );
NAND3X1 NAND3X1_2790 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf1_), .B(_12293_), .C(_12295_), .Y(_12305_) );
NAND3X1 NAND3X1_2791 ( .gnd(gnd), .vdd(vdd), .A(_12086_), .B(_12305_), .C(_12304_), .Y(_12306_) );
AOI21X1 AOI21X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_12306_), .B(_12303_), .C(_12277_), .Y(_12307_) );
INVX2 INVX2_412 ( .gnd(gnd), .vdd(vdd), .A(_12307_), .Y(_12308_) );
NAND3X1 NAND3X1_2792 ( .gnd(gnd), .vdd(vdd), .A(_12277_), .B(_12306_), .C(_12303_), .Y(_12309_) );
AOI21X1 AOI21X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_12309_), .B(_12308_), .C(bloque_datos_19_bF_buf3_), .Y(_12310_) );
INVX1 INVX1_1706 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf2_), .Y(_12311_) );
INVX2 INVX2_413 ( .gnd(gnd), .vdd(vdd), .A(_12309_), .Y(_12312_) );
NOR3X1 NOR3X1_362 ( .gnd(gnd), .vdd(vdd), .A(_12311_), .B(_12307_), .C(_12312_), .Y(_12313_) );
OAI21X1 OAI21X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_12313_), .B(_12310_), .C(_12100_), .Y(_12314_) );
OAI21X1 OAI21X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_12312_), .B(_12307_), .C(_12311_), .Y(_12315_) );
NAND3X1 NAND3X1_2793 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf1_), .B(_12309_), .C(_12308_), .Y(_12316_) );
NAND3X1 NAND3X1_2794 ( .gnd(gnd), .vdd(vdd), .A(_12104_), .B(_12315_), .C(_12316_), .Y(_12317_) );
AOI21X1 AOI21X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_12317_), .B(_12314_), .C(_12276_), .Y(_12318_) );
NAND2X1 NAND2X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_12317_), .B(_12314_), .Y(_12319_) );
NOR2X1 NOR2X1_934 ( .gnd(gnd), .vdd(vdd), .A(_12275_), .B(_12319_), .Y(_12320_) );
OAI21X1 OAI21X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_12320_), .B(_12318_), .C(bloque_datos_35_bF_buf2_), .Y(_12321_) );
INVX1 INVX1_1707 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf1_), .Y(_12322_) );
INVX1 INVX1_1708 ( .gnd(gnd), .vdd(vdd), .A(_12314_), .Y(_12323_) );
INVX1 INVX1_1709 ( .gnd(gnd), .vdd(vdd), .A(_12317_), .Y(_12324_) );
OAI21X1 OAI21X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_12323_), .B(_12324_), .C(_12275_), .Y(_12325_) );
NAND3X1 NAND3X1_2795 ( .gnd(gnd), .vdd(vdd), .A(_12317_), .B(_12314_), .C(_12276_), .Y(_12326_) );
NAND3X1 NAND3X1_2796 ( .gnd(gnd), .vdd(vdd), .A(_12322_), .B(_12326_), .C(_12325_), .Y(_12327_) );
NAND3X1 NAND3X1_2797 ( .gnd(gnd), .vdd(vdd), .A(_12116_), .B(_12327_), .C(_12321_), .Y(_12328_) );
OAI21X1 OAI21X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_12320_), .B(_12318_), .C(_12322_), .Y(_12329_) );
NAND3X1 NAND3X1_2798 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf0_), .B(_12326_), .C(_12325_), .Y(_12330_) );
NAND3X1 NAND3X1_2799 ( .gnd(gnd), .vdd(vdd), .A(_12113_), .B(_12330_), .C(_12329_), .Y(_12331_) );
NAND2X1 NAND2X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_12328_), .B(_12331_), .Y(_12332_) );
NAND2X1 NAND2X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_12332_), .B(_12274_), .Y(_12333_) );
OR2X2 OR2X2_282 ( .gnd(gnd), .vdd(vdd), .A(_12274_), .B(_12332_), .Y(_12334_) );
NAND2X1 NAND2X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_12333_), .B(_12334_), .Y(_12335_) );
XNOR2X1 XNOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_12335_), .B(bloque_datos_51_bF_buf2_), .Y(_12336_) );
OR2X2 OR2X2_283 ( .gnd(gnd), .vdd(vdd), .A(_12336_), .B(_12273_), .Y(_12337_) );
NOR2X1 NOR2X1_935 ( .gnd(gnd), .vdd(vdd), .A(_12119_), .B(_12123_), .Y(_12338_) );
INVX2 INVX2_414 ( .gnd(gnd), .vdd(vdd), .A(_12338_), .Y(_12339_) );
OAI21X1 OAI21X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_12122_), .B(_12339_), .C(_12336_), .Y(_12340_) );
AOI21X1 AOI21X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_12340_), .B(_12337_), .C(_12272_), .Y(_12341_) );
INVX2 INVX2_415 ( .gnd(gnd), .vdd(vdd), .A(_12272_), .Y(_12342_) );
NOR2X1 NOR2X1_936 ( .gnd(gnd), .vdd(vdd), .A(_12273_), .B(_12336_), .Y(_12343_) );
NAND2X1 NAND2X1_1616 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf1_), .B(_12335_), .Y(_12344_) );
OR2X2 OR2X2_284 ( .gnd(gnd), .vdd(vdd), .A(_12335_), .B(bloque_datos_51_bF_buf0_), .Y(_12345_) );
AOI21X1 AOI21X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_12344_), .B(_12345_), .C(_12124_), .Y(_12346_) );
NOR3X1 NOR3X1_363 ( .gnd(gnd), .vdd(vdd), .A(_12342_), .B(_12346_), .C(_12343_), .Y(_12347_) );
OAI21X1 OAI21X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_12341_), .B(_12347_), .C(bloque_datos_67_bF_buf0_), .Y(_12348_) );
INVX1 INVX1_1710 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf4_), .Y(_12349_) );
NOR2X1 NOR2X1_937 ( .gnd(gnd), .vdd(vdd), .A(_12347_), .B(_12341_), .Y(_12350_) );
NAND2X1 NAND2X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_12349_), .B(_12350_), .Y(_12351_) );
NAND3X1 NAND3X1_2800 ( .gnd(gnd), .vdd(vdd), .A(_12140_), .B(_12348_), .C(_12351_), .Y(_12352_) );
OAI21X1 OAI21X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_12341_), .B(_12347_), .C(_12349_), .Y(_12353_) );
NAND2X1 NAND2X1_1618 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf3_), .B(_12350_), .Y(_12354_) );
NAND3X1 NAND3X1_2801 ( .gnd(gnd), .vdd(vdd), .A(_12136_), .B(_12353_), .C(_12354_), .Y(_12355_) );
AOI21X1 AOI21X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_12355_), .B(_12352_), .C(_12271_), .Y(_12356_) );
NAND3X1 NAND3X1_2802 ( .gnd(gnd), .vdd(vdd), .A(_12271_), .B(_12355_), .C(_12352_), .Y(_12357_) );
INVX2 INVX2_416 ( .gnd(gnd), .vdd(vdd), .A(_12357_), .Y(_12358_) );
OAI21X1 OAI21X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_12358_), .B(_12356_), .C(bloque_datos_83_bF_buf1_), .Y(_12359_) );
INVX1 INVX1_1711 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf0_), .Y(_12360_) );
INVX2 INVX2_417 ( .gnd(gnd), .vdd(vdd), .A(_12356_), .Y(_12361_) );
NAND3X1 NAND3X1_2803 ( .gnd(gnd), .vdd(vdd), .A(_12360_), .B(_12357_), .C(_12361_), .Y(_12362_) );
NAND3X1 NAND3X1_2804 ( .gnd(gnd), .vdd(vdd), .A(_12151_), .B(_12362_), .C(_12359_), .Y(_12363_) );
INVX1 INVX1_1712 ( .gnd(gnd), .vdd(vdd), .A(_12151_), .Y(_12364_) );
OAI21X1 OAI21X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_12358_), .B(_12356_), .C(_12360_), .Y(_12365_) );
NAND3X1 NAND3X1_2805 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf5_), .B(_12357_), .C(_12361_), .Y(_12366_) );
NAND3X1 NAND3X1_2806 ( .gnd(gnd), .vdd(vdd), .A(_12364_), .B(_12366_), .C(_12365_), .Y(_12367_) );
AOI21X1 AOI21X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_12363_), .B(_12367_), .C(_12270_), .Y(_12368_) );
NAND3X1 NAND3X1_2807 ( .gnd(gnd), .vdd(vdd), .A(_12270_), .B(_12363_), .C(_12367_), .Y(_12369_) );
INVX2 INVX2_418 ( .gnd(gnd), .vdd(vdd), .A(_12369_), .Y(_12370_) );
OAI21X1 OAI21X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_12370_), .B(_12368_), .C(_12269_), .Y(_12371_) );
INVX1 INVX1_1713 ( .gnd(gnd), .vdd(vdd), .A(_12368_), .Y(_12372_) );
NAND3X1 NAND3X1_2808 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_131_), .B(_12369_), .C(_12372_), .Y(_12373_) );
NAND2X1 NAND2X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_12373_), .B(_12371_), .Y(_12374_) );
NAND2X1 NAND2X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_12163_), .B(_12374_), .Y(_12375_) );
INVX1 INVX1_1714 ( .gnd(gnd), .vdd(vdd), .A(_12163_), .Y(_12376_) );
NAND3X1 NAND3X1_2809 ( .gnd(gnd), .vdd(vdd), .A(_12376_), .B(_12373_), .C(_12371_), .Y(_12377_) );
NAND3X1 NAND3X1_2810 ( .gnd(gnd), .vdd(vdd), .A(_12377_), .B(_12375_), .C(_12268_), .Y(_12378_) );
INVX1 INVX1_1715 ( .gnd(gnd), .vdd(vdd), .A(_12378_), .Y(_12379_) );
AND2X2 AND2X2_272 ( .gnd(gnd), .vdd(vdd), .A(_12375_), .B(_12377_), .Y(_12380_) );
NOR2X1 NOR2X1_938 ( .gnd(gnd), .vdd(vdd), .A(_12268_), .B(_12380_), .Y(_12381_) );
OAI21X1 OAI21X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_12381_), .B(_12379_), .C(_12267_), .Y(_12382_) );
NOR3X1 NOR3X1_364 ( .gnd(gnd), .vdd(vdd), .A(_12267_), .B(_12379_), .C(_12381_), .Y(_12383_) );
INVX2 INVX2_419 ( .gnd(gnd), .vdd(vdd), .A(_12383_), .Y(_12384_) );
NAND3X1 NAND3X1_2811 ( .gnd(gnd), .vdd(vdd), .A(_12175_), .B(_12382_), .C(_12384_), .Y(_12385_) );
INVX1 INVX1_1716 ( .gnd(gnd), .vdd(vdd), .A(_12175_), .Y(_12386_) );
INVX1 INVX1_1717 ( .gnd(gnd), .vdd(vdd), .A(_12382_), .Y(_12387_) );
OAI21X1 OAI21X1_1958 ( .gnd(gnd), .vdd(vdd), .A(_12387_), .B(_12383_), .C(_12386_), .Y(_12388_) );
NAND3X1 NAND3X1_2812 ( .gnd(gnd), .vdd(vdd), .A(_12388_), .B(_12266_), .C(_12385_), .Y(_12389_) );
INVX1 INVX1_1718 ( .gnd(gnd), .vdd(vdd), .A(_12389_), .Y(_12390_) );
AOI21X1 AOI21X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_12388_), .B(_12385_), .C(_12266_), .Y(_12391_) );
OAI21X1 OAI21X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_12390_), .B(_12391_), .C(_12264_), .Y(_12392_) );
NOR2X1 NOR2X1_939 ( .gnd(gnd), .vdd(vdd), .A(_12391_), .B(_12390_), .Y(_12393_) );
NAND2X1 NAND2X1_1621 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_163_), .B(_12393_), .Y(_12394_) );
NAND2X1 NAND2X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_12392_), .B(_12394_), .Y(_12395_) );
NOR2X1 NOR2X1_940 ( .gnd(gnd), .vdd(vdd), .A(_12185_), .B(_12395_), .Y(_12396_) );
INVX2 INVX2_420 ( .gnd(gnd), .vdd(vdd), .A(_12184_), .Y(_12397_) );
OAI21X1 OAI21X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_12057_), .B(_12397_), .C(_12395_), .Y(_12398_) );
INVX2 INVX2_421 ( .gnd(gnd), .vdd(vdd), .A(_12398_), .Y(_12399_) );
NOR2X1 NOR2X1_941 ( .gnd(gnd), .vdd(vdd), .A(_12396_), .B(_12399_), .Y(_12400_) );
OAI21X1 OAI21X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_12191_), .B(_12263_), .C(_12400_), .Y(_12401_) );
AOI21X1 AOI21X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_12016_), .B(_12189_), .C(_12263_), .Y(_12402_) );
OAI21X1 OAI21X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_12399_), .B(_12396_), .C(_12402_), .Y(_12403_) );
NAND2X1 NAND2X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_12403_), .B(_12401_), .Y(_12404_) );
NAND2X1 NAND2X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_12262_), .B(_12404_), .Y(_12405_) );
NOR2X1 NOR2X1_942 ( .gnd(gnd), .vdd(vdd), .A(_12262_), .B(_12404_), .Y(_12406_) );
INVX2 INVX2_422 ( .gnd(gnd), .vdd(vdd), .A(_12406_), .Y(_12407_) );
NAND3X1 NAND3X1_2813 ( .gnd(gnd), .vdd(vdd), .A(_12198_), .B(_12405_), .C(_12407_), .Y(_12408_) );
INVX1 INVX1_1719 ( .gnd(gnd), .vdd(vdd), .A(_12405_), .Y(_12409_) );
OAI21X1 OAI21X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_12409_), .B(_12406_), .C(_12195_), .Y(_12410_) );
NAND2X1 NAND2X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_12410_), .B(_12408_), .Y(_12411_) );
NOR2X1 NOR2X1_943 ( .gnd(gnd), .vdd(vdd), .A(_12261_), .B(_12411_), .Y(_12412_) );
INVX1 INVX1_1720 ( .gnd(gnd), .vdd(vdd), .A(_12408_), .Y(_12413_) );
INVX1 INVX1_1721 ( .gnd(gnd), .vdd(vdd), .A(_12410_), .Y(_12414_) );
OAI21X1 OAI21X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_12413_), .B(_12414_), .C(_12261_), .Y(_12415_) );
INVX1 INVX1_1722 ( .gnd(gnd), .vdd(vdd), .A(_12415_), .Y(_12416_) );
OAI21X1 OAI21X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_12416_), .B(_12412_), .C(_12260_), .Y(_12417_) );
NOR2X1 NOR2X1_944 ( .gnd(gnd), .vdd(vdd), .A(_12412_), .B(_12416_), .Y(_12418_) );
NAND2X1 NAND2X1_1626 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_195_), .B(_12418_), .Y(_12419_) );
NAND2X1 NAND2X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_12417_), .B(_12419_), .Y(_12420_) );
OR2X2 OR2X2_285 ( .gnd(gnd), .vdd(vdd), .A(_12420_), .B(_12259_), .Y(_12421_) );
AOI21X1 AOI21X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_12417_), .B(_12419_), .C(_12205_), .Y(_12422_) );
INVX1 INVX1_1723 ( .gnd(gnd), .vdd(vdd), .A(_12422_), .Y(_12423_) );
NAND2X1 NAND2X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_12423_), .B(_12421_), .Y(_12424_) );
NOR2X1 NOR2X1_945 ( .gnd(gnd), .vdd(vdd), .A(_12258_), .B(_12424_), .Y(_12425_) );
NOR2X1 NOR2X1_946 ( .gnd(gnd), .vdd(vdd), .A(_12259_), .B(_12420_), .Y(_12426_) );
OAI21X1 OAI21X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_12426_), .B(_12422_), .C(_12258_), .Y(_12427_) );
INVX2 INVX2_423 ( .gnd(gnd), .vdd(vdd), .A(_12427_), .Y(_12428_) );
OAI21X1 OAI21X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_12425_), .B(_12428_), .C(_12256_), .Y(_12429_) );
INVX1 INVX1_1724 ( .gnd(gnd), .vdd(vdd), .A(_12429_), .Y(_12430_) );
NOR2X1 NOR2X1_947 ( .gnd(gnd), .vdd(vdd), .A(_12422_), .B(_12426_), .Y(_12431_) );
OAI21X1 OAI21X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_12257_), .B(_12210_), .C(_12431_), .Y(_12432_) );
NAND2X1 NAND2X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_12427_), .B(_12432_), .Y(_12433_) );
NOR2X1 NOR2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_12256_), .B(_12433_), .Y(_12434_) );
NOR3X1 NOR3X1_365 ( .gnd(gnd), .vdd(vdd), .A(_12255_), .B(_12434_), .C(_12430_), .Y(_12435_) );
NOR2X1 NOR2X1_949 ( .gnd(gnd), .vdd(vdd), .A(_12428_), .B(_12425_), .Y(_12436_) );
NAND2X1 NAND2X1_1630 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_211_), .B(_12436_), .Y(_12437_) );
AOI21X1 AOI21X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_12429_), .B(_12437_), .C(_12215_), .Y(_12438_) );
NOR2X1 NOR2X1_950 ( .gnd(gnd), .vdd(vdd), .A(_12438_), .B(_12435_), .Y(_12439_) );
AND2X2 AND2X2_273 ( .gnd(gnd), .vdd(vdd), .A(_12439_), .B(_12254_), .Y(_12440_) );
INVX1 INVX1_1725 ( .gnd(gnd), .vdd(vdd), .A(_12254_), .Y(_12441_) );
OAI21X1 OAI21X1_1969 ( .gnd(gnd), .vdd(vdd), .A(_12435_), .B(_12438_), .C(_12441_), .Y(_12442_) );
INVX2 INVX2_424 ( .gnd(gnd), .vdd(vdd), .A(_12442_), .Y(_12443_) );
OAI21X1 OAI21X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_12440_), .B(_12443_), .C(_12253_), .Y(_12444_) );
NOR2X1 NOR2X1_951 ( .gnd(gnd), .vdd(vdd), .A(_12443_), .B(_12440_), .Y(_12445_) );
NAND2X1 NAND2X1_1631 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_227_), .B(_12445_), .Y(_12446_) );
NAND3X1 NAND3X1_2814 ( .gnd(gnd), .vdd(vdd), .A(_12228_), .B(_12444_), .C(_12446_), .Y(_12447_) );
NAND2X1 NAND2X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_12444_), .B(_12446_), .Y(_12448_) );
NAND2X1 NAND2X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_12226_), .B(_12448_), .Y(_12449_) );
NAND3X1 NAND3X1_2815 ( .gnd(gnd), .vdd(vdd), .A(_12252_), .B(_12447_), .C(_12449_), .Y(_12450_) );
INVX2 INVX2_425 ( .gnd(gnd), .vdd(vdd), .A(_12450_), .Y(_12451_) );
AND2X2 AND2X2_274 ( .gnd(gnd), .vdd(vdd), .A(_12230_), .B(_12227_), .Y(_12452_) );
INVX1 INVX1_1726 ( .gnd(gnd), .vdd(vdd), .A(_12447_), .Y(_12453_) );
AOI21X1 AOI21X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_12444_), .B(_12446_), .C(_12228_), .Y(_12454_) );
OAI21X1 OAI21X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_12453_), .B(_12454_), .C(_12452_), .Y(_12455_) );
INVX2 INVX2_426 ( .gnd(gnd), .vdd(vdd), .A(_12455_), .Y(_12456_) );
OAI21X1 OAI21X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_12456_), .B(_12451_), .C(_12251_), .Y(_12457_) );
NOR2X1 NOR2X1_952 ( .gnd(gnd), .vdd(vdd), .A(_12451_), .B(_12456_), .Y(_12458_) );
NAND2X1 NAND2X1_1634 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_243_), .B(_12458_), .Y(_12459_) );
NAND2X1 NAND2X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_12457_), .B(_12459_), .Y(_12460_) );
OR2X2 OR2X2_286 ( .gnd(gnd), .vdd(vdd), .A(_12460_), .B(_12235_), .Y(_12461_) );
INVX2 INVX2_427 ( .gnd(gnd), .vdd(vdd), .A(_12234_), .Y(_12462_) );
OAI21X1 OAI21X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_12462_), .B(_12054_), .C(_12460_), .Y(_12463_) );
AOI21X1 AOI21X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_12463_), .B(_12461_), .C(_12250_), .Y(_12464_) );
INVX1 INVX1_1727 ( .gnd(gnd), .vdd(vdd), .A(_12250_), .Y(_12465_) );
NAND2X1 NAND2X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_12463_), .B(_12461_), .Y(_12466_) );
NOR2X1 NOR2X1_953 ( .gnd(gnd), .vdd(vdd), .A(_12465_), .B(_12466_), .Y(_12467_) );
NOR2X1 NOR2X1_954 ( .gnd(gnd), .vdd(vdd), .A(_12464_), .B(_12467_), .Y(_12468_) );
INVX2 INVX2_428 ( .gnd(gnd), .vdd(vdd), .A(_12468_), .Y(module_2_H_15_) );
NOR2X1 NOR2X1_955 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_240_), .B(_12240_), .Y(_12469_) );
OAI21X1 OAI21X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_12242_), .B(_12053_), .C(_12469_), .Y(_12470_) );
NAND2X1 NAND2X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_12470_), .B(_12244_), .Y(_12471_) );
INVX2 INVX2_429 ( .gnd(gnd), .vdd(vdd), .A(_12471_), .Y(module_2_H_13_) );
NAND2X1 NAND2X1_1638 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_240_), .B(_12240_), .Y(_12472_) );
INVX1 INVX1_1728 ( .gnd(gnd), .vdd(vdd), .A(_12472_), .Y(_12473_) );
NOR2X1 NOR2X1_956 ( .gnd(gnd), .vdd(vdd), .A(_12469_), .B(_12473_), .Y(module_2_H_0_) );
INVX1 INVX1_1729 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_0_), .Y(module_2_H_12_) );
INVX1 INVX1_1730 ( .gnd(gnd), .vdd(vdd), .A(_12244_), .Y(_12474_) );
OAI21X1 OAI21X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_12469_), .B(_12473_), .C(module_2_H_13_), .Y(_12475_) );
INVX2 INVX2_430 ( .gnd(gnd), .vdd(vdd), .A(_12475_), .Y(_12476_) );
AOI21X1 AOI21X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_12474_), .B(_12472_), .C(_12476_), .Y(module_2_H_1_) );
NAND3X1 NAND3X1_2816 ( .gnd(gnd), .vdd(vdd), .A(_12236_), .B(_12474_), .C(_12248_), .Y(_12477_) );
INVX1 INVX1_1731 ( .gnd(gnd), .vdd(vdd), .A(_12236_), .Y(_12478_) );
OAI21X1 OAI21X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_12249_), .B(_12478_), .C(_12244_), .Y(_12479_) );
AND2X2 AND2X2_275 ( .gnd(gnd), .vdd(vdd), .A(_12479_), .B(_12477_), .Y(module_2_H_14_) );
NAND2X1 NAND2X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_12476_), .B(module_2_H_14_), .Y(_12480_) );
INVX1 INVX1_1732 ( .gnd(gnd), .vdd(vdd), .A(_12480_), .Y(_12481_) );
NOR2X1 NOR2X1_957 ( .gnd(gnd), .vdd(vdd), .A(_12476_), .B(module_2_H_14_), .Y(_12482_) );
NOR2X1 NOR2X1_958 ( .gnd(gnd), .vdd(vdd), .A(_12482_), .B(_12481_), .Y(module_2_H_2_) );
NOR3X1 NOR3X1_366 ( .gnd(gnd), .vdd(vdd), .A(_12480_), .B(_12464_), .C(_12467_), .Y(_12483_) );
NOR2X1 NOR2X1_959 ( .gnd(gnd), .vdd(vdd), .A(_12481_), .B(_12468_), .Y(_12484_) );
NOR2X1 NOR2X1_960 ( .gnd(gnd), .vdd(vdd), .A(_12483_), .B(_12484_), .Y(module_2_H_3_) );
AOI21X1 AOI21X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_12457_), .B(_12459_), .C(_12247_), .Y(_12485_) );
OAI21X1 OAI21X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_12465_), .B(_12485_), .C(_12461_), .Y(_12486_) );
INVX1 INVX1_1733 ( .gnd(gnd), .vdd(vdd), .A(_12459_), .Y(_12487_) );
AOI21X1 AOI21X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_12252_), .B(_12449_), .C(_12453_), .Y(_12488_) );
OAI21X1 OAI21X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_12430_), .B(_12434_), .C(_12255_), .Y(_12489_) );
AOI21X1 AOI21X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_12254_), .B(_12489_), .C(_12435_), .Y(_12490_) );
INVX1 INVX1_1734 ( .gnd(gnd), .vdd(vdd), .A(_12258_), .Y(_12491_) );
AOI21X1 AOI21X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_12491_), .B(_12423_), .C(_12426_), .Y(_12492_) );
NAND2X1 NAND2X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_12196_), .B(_12200_), .Y(_12493_) );
AOI21X1 AOI21X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_12493_), .B(_12410_), .C(_12413_), .Y(_12494_) );
INVX1 INVX1_1735 ( .gnd(gnd), .vdd(vdd), .A(_12396_), .Y(_12495_) );
OAI21X1 OAI21X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_12399_), .B(_12402_), .C(_12495_), .Y(_12496_) );
INVX1 INVX1_1736 ( .gnd(gnd), .vdd(vdd), .A(_12496_), .Y(_12497_) );
AND2X2 AND2X2_276 ( .gnd(gnd), .vdd(vdd), .A(_12389_), .B(_12385_), .Y(_12498_) );
NAND2X1 NAND2X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_12375_), .B(_12378_), .Y(_12499_) );
AND2X2 AND2X2_277 ( .gnd(gnd), .vdd(vdd), .A(_12369_), .B(_12363_), .Y(_12500_) );
INVX2 INVX2_431 ( .gnd(gnd), .vdd(vdd), .A(_12365_), .Y(_12501_) );
AOI21X1 AOI21X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_12353_), .B(_12354_), .C(_12136_), .Y(_12502_) );
AOI21X1 AOI21X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_12271_), .B(_12355_), .C(_12502_), .Y(_12503_) );
INVX2 INVX2_432 ( .gnd(gnd), .vdd(vdd), .A(_12353_), .Y(_12504_) );
AOI21X1 AOI21X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_12272_), .B(_12340_), .C(_12343_), .Y(_12505_) );
INVX1 INVX1_1737 ( .gnd(gnd), .vdd(vdd), .A(_12335_), .Y(_12506_) );
NOR2X1 NOR2X1_961 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf4_), .B(_12506_), .Y(_12507_) );
NAND2X1 NAND2X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_12114_), .B(_12118_), .Y(_12508_) );
INVX1 INVX1_1738 ( .gnd(gnd), .vdd(vdd), .A(_12328_), .Y(_12509_) );
AOI21X1 AOI21X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_12331_), .B(_12508_), .C(_12509_), .Y(_12510_) );
INVX2 INVX2_433 ( .gnd(gnd), .vdd(vdd), .A(_12329_), .Y(_12511_) );
AOI21X1 AOI21X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_12317_), .B(_12276_), .C(_12323_), .Y(_12512_) );
AOI21X1 AOI21X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_12305_), .B(_12304_), .C(_12086_), .Y(_12513_) );
AOI21X1 AOI21X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_12306_), .B(_12277_), .C(_12513_), .Y(_12514_) );
OAI21X1 OAI21X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_12290_), .B(_12291_), .C(_12077_), .Y(_12515_) );
OAI21X1 OAI21X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_12279_), .B(_12292_), .C(_12515_), .Y(_12516_) );
INVX1 INVX1_1739 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_4_), .Y(_12517_) );
OAI21X1 OAI21X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_12069_), .B(_12281_), .C(_12517_), .Y(_12518_) );
NAND2X1 NAND2X1_1643 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_4_), .B(_12282_), .Y(_12519_) );
AOI21X1 AOI21X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_12518_), .B(_12519_), .C(_11312_), .Y(_12520_) );
INVX1 INVX1_1740 ( .gnd(gnd), .vdd(vdd), .A(_12518_), .Y(_12521_) );
NOR3X1 NOR3X1_367 ( .gnd(gnd), .vdd(vdd), .A(_12281_), .B(_12517_), .C(_12069_), .Y(_12522_) );
NOR3X1 NOR3X1_368 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_0_), .B(_12522_), .C(_12521_), .Y(_12523_) );
OAI21X1 OAI21X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_12523_), .B(_12520_), .C(module_2_W_20_), .Y(_12524_) );
INVX1 INVX1_1741 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_20_), .Y(_12525_) );
OAI21X1 OAI21X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_12521_), .B(_12522_), .C(module_2_W_0_), .Y(_12526_) );
NAND3X1 NAND3X1_2817 ( .gnd(gnd), .vdd(vdd), .A(_11312_), .B(_12518_), .C(_12519_), .Y(_12527_) );
NAND3X1 NAND3X1_2818 ( .gnd(gnd), .vdd(vdd), .A(_12525_), .B(_12527_), .C(_12526_), .Y(_12528_) );
NAND3X1 NAND3X1_2819 ( .gnd(gnd), .vdd(vdd), .A(_12284_), .B(_12528_), .C(_12524_), .Y(_12529_) );
OAI21X1 OAI21X1_1985 ( .gnd(gnd), .vdd(vdd), .A(_12523_), .B(_12520_), .C(_12525_), .Y(_12530_) );
NAND3X1 NAND3X1_2820 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_20_), .B(_12527_), .C(_12526_), .Y(_12531_) );
NAND3X1 NAND3X1_2821 ( .gnd(gnd), .vdd(vdd), .A(_12290_), .B(_12531_), .C(_12530_), .Y(_12532_) );
NAND3X1 NAND3X1_2822 ( .gnd(gnd), .vdd(vdd), .A(_12529_), .B(_12532_), .C(_12516_), .Y(_12533_) );
NAND3X1 NAND3X1_2823 ( .gnd(gnd), .vdd(vdd), .A(_12074_), .B(_12284_), .C(_12286_), .Y(_12534_) );
AOI21X1 AOI21X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_12534_), .B(_12300_), .C(_12287_), .Y(_12535_) );
NAND3X1 NAND3X1_2824 ( .gnd(gnd), .vdd(vdd), .A(_12290_), .B(_12528_), .C(_12524_), .Y(_12536_) );
NAND3X1 NAND3X1_2825 ( .gnd(gnd), .vdd(vdd), .A(_12284_), .B(_12531_), .C(_12530_), .Y(_12537_) );
NAND3X1 NAND3X1_2826 ( .gnd(gnd), .vdd(vdd), .A(_12535_), .B(_12536_), .C(_12537_), .Y(_12538_) );
XNOR2X1 XNOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_10614_), .B(module_2_W_8_), .Y(_12539_) );
INVX1 INVX1_1742 ( .gnd(gnd), .vdd(vdd), .A(_12539_), .Y(_12540_) );
NAND3X1 NAND3X1_2827 ( .gnd(gnd), .vdd(vdd), .A(_12540_), .B(_12538_), .C(_12533_), .Y(_12541_) );
AOI21X1 AOI21X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_12536_), .B(_12537_), .C(_12535_), .Y(_12542_) );
AOI21X1 AOI21X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_12529_), .B(_12532_), .C(_12516_), .Y(_12543_) );
OAI21X1 OAI21X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_12542_), .B(_12543_), .C(_12539_), .Y(_12544_) );
AOI21X1 AOI21X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_12541_), .B(_12544_), .C(bloque_datos_4_bF_buf3_), .Y(_12545_) );
INVX1 INVX1_1743 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf2_), .Y(_12546_) );
NAND3X1 NAND3X1_2828 ( .gnd(gnd), .vdd(vdd), .A(_12539_), .B(_12538_), .C(_12533_), .Y(_12547_) );
OAI21X1 OAI21X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_12542_), .B(_12543_), .C(_12540_), .Y(_12548_) );
AOI21X1 AOI21X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_12547_), .B(_12548_), .C(_12546_), .Y(_12549_) );
OAI21X1 OAI21X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_12545_), .B(_12549_), .C(_12296_), .Y(_12550_) );
NAND3X1 NAND3X1_2829 ( .gnd(gnd), .vdd(vdd), .A(_12546_), .B(_12547_), .C(_12548_), .Y(_12551_) );
NAND3X1 NAND3X1_2830 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf1_), .B(_12541_), .C(_12544_), .Y(_12552_) );
NAND3X1 NAND3X1_2831 ( .gnd(gnd), .vdd(vdd), .A(_12304_), .B(_12551_), .C(_12552_), .Y(_12553_) );
NAND3X1 NAND3X1_2832 ( .gnd(gnd), .vdd(vdd), .A(_12514_), .B(_12553_), .C(_12550_), .Y(_12554_) );
AOI21X1 AOI21X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_12090_), .B(_12065_), .C(_12097_), .Y(_12555_) );
NOR3X1 NOR3X1_369 ( .gnd(gnd), .vdd(vdd), .A(_12089_), .B(_12296_), .C(_12302_), .Y(_12556_) );
OAI21X1 OAI21X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_12556_), .B(_12555_), .C(_12303_), .Y(_12557_) );
OAI21X1 OAI21X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_12545_), .B(_12549_), .C(_12304_), .Y(_12558_) );
NAND3X1 NAND3X1_2833 ( .gnd(gnd), .vdd(vdd), .A(_12296_), .B(_12551_), .C(_12552_), .Y(_12559_) );
NAND3X1 NAND3X1_2834 ( .gnd(gnd), .vdd(vdd), .A(_12559_), .B(_12558_), .C(_12557_), .Y(_12560_) );
NOR2X1 NOR2X1_962 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_24_), .B(module_2_W_8_), .Y(_12561_) );
INVX1 INVX1_1744 ( .gnd(gnd), .vdd(vdd), .A(_12561_), .Y(_12562_) );
NAND2X1 NAND2X1_1644 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_24_), .B(module_2_W_8_), .Y(_12563_) );
NAND2X1 NAND2X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_12563_), .B(_12562_), .Y(_12564_) );
XNOR2X1 XNOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_10636_), .B(_12564_), .Y(_12565_) );
NAND3X1 NAND3X1_2835 ( .gnd(gnd), .vdd(vdd), .A(_12565_), .B(_12554_), .C(_12560_), .Y(_12566_) );
AOI21X1 AOI21X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_12559_), .B(_12558_), .C(_12557_), .Y(_12567_) );
AOI21X1 AOI21X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_12553_), .B(_12550_), .C(_12514_), .Y(_12568_) );
INVX1 INVX1_1745 ( .gnd(gnd), .vdd(vdd), .A(_12565_), .Y(_12569_) );
OAI21X1 OAI21X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_12567_), .B(_12568_), .C(_12569_), .Y(_12570_) );
AOI21X1 AOI21X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_12566_), .B(_12570_), .C(bloque_datos_20_bF_buf3_), .Y(_12571_) );
INVX1 INVX1_1746 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf2_), .Y(_12572_) );
OAI21X1 OAI21X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_12567_), .B(_12568_), .C(_12565_), .Y(_12573_) );
NAND3X1 NAND3X1_2836 ( .gnd(gnd), .vdd(vdd), .A(_12569_), .B(_12554_), .C(_12560_), .Y(_12574_) );
AOI21X1 AOI21X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_12574_), .B(_12573_), .C(_12572_), .Y(_12575_) );
OAI21X1 OAI21X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_12571_), .B(_12575_), .C(_12310_), .Y(_12576_) );
NAND3X1 NAND3X1_2837 ( .gnd(gnd), .vdd(vdd), .A(_12572_), .B(_12574_), .C(_12573_), .Y(_12577_) );
NAND3X1 NAND3X1_2838 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf1_), .B(_12566_), .C(_12570_), .Y(_12578_) );
NAND3X1 NAND3X1_2839 ( .gnd(gnd), .vdd(vdd), .A(_12315_), .B(_12577_), .C(_12578_), .Y(_12579_) );
NAND3X1 NAND3X1_2840 ( .gnd(gnd), .vdd(vdd), .A(_12579_), .B(_12576_), .C(_12512_), .Y(_12580_) );
OAI21X1 OAI21X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_12324_), .B(_12275_), .C(_12314_), .Y(_12581_) );
OAI21X1 OAI21X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_12571_), .B(_12575_), .C(_12315_), .Y(_12582_) );
NAND3X1 NAND3X1_2841 ( .gnd(gnd), .vdd(vdd), .A(_12310_), .B(_12577_), .C(_12578_), .Y(_12583_) );
NAND3X1 NAND3X1_2842 ( .gnd(gnd), .vdd(vdd), .A(_12583_), .B(_12581_), .C(_12582_), .Y(_12584_) );
INVX1 INVX1_1747 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .Y(_12585_) );
OR2X2 OR2X2_287 ( .gnd(gnd), .vdd(vdd), .A(_12564_), .B(_12585_), .Y(_12586_) );
NAND2X1 NAND2X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_12585_), .B(_12564_), .Y(_12587_) );
NAND2X1 NAND2X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_12587_), .B(_12586_), .Y(_12588_) );
INVX2 INVX2_434 ( .gnd(gnd), .vdd(vdd), .A(_12588_), .Y(_12589_) );
XNOR2X1 XNOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_10667_), .B(_12589_), .Y(_12590_) );
NAND3X1 NAND3X1_2843 ( .gnd(gnd), .vdd(vdd), .A(_12590_), .B(_12584_), .C(_12580_), .Y(_12591_) );
AOI21X1 AOI21X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_12583_), .B(_12582_), .C(_12581_), .Y(_8782_) );
AOI21X1 AOI21X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_12579_), .B(_12576_), .C(_12512_), .Y(_8783_) );
INVX1 INVX1_1748 ( .gnd(gnd), .vdd(vdd), .A(_12590_), .Y(_8784_) );
OAI21X1 OAI21X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_8782_), .B(_8783_), .C(_8784_), .Y(_8785_) );
AOI21X1 AOI21X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_12591_), .B(_8785_), .C(bloque_datos_36_bF_buf1_), .Y(_8786_) );
INVX1 INVX1_1749 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf0_), .Y(_8787_) );
NAND3X1 NAND3X1_2844 ( .gnd(gnd), .vdd(vdd), .A(_8784_), .B(_12584_), .C(_12580_), .Y(_8788_) );
OAI21X1 OAI21X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_8782_), .B(_8783_), .C(_12590_), .Y(_8789_) );
AOI21X1 AOI21X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_8788_), .B(_8789_), .C(_8787_), .Y(_8790_) );
OAI21X1 OAI21X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_8786_), .B(_8790_), .C(_12511_), .Y(_8791_) );
NAND3X1 NAND3X1_2845 ( .gnd(gnd), .vdd(vdd), .A(_8787_), .B(_8788_), .C(_8789_), .Y(_8792_) );
NAND3X1 NAND3X1_2846 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf3_), .B(_12591_), .C(_8785_), .Y(_8793_) );
NAND3X1 NAND3X1_2847 ( .gnd(gnd), .vdd(vdd), .A(_12329_), .B(_8792_), .C(_8793_), .Y(_8794_) );
NAND3X1 NAND3X1_2848 ( .gnd(gnd), .vdd(vdd), .A(_12510_), .B(_8794_), .C(_8791_), .Y(_8795_) );
OAI21X1 OAI21X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_12274_), .B(_12332_), .C(_12328_), .Y(_8796_) );
OAI21X1 OAI21X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_8786_), .B(_8790_), .C(_12329_), .Y(_8797_) );
NAND3X1 NAND3X1_2849 ( .gnd(gnd), .vdd(vdd), .A(_12511_), .B(_8792_), .C(_8793_), .Y(_8798_) );
NAND3X1 NAND3X1_2850 ( .gnd(gnd), .vdd(vdd), .A(_8796_), .B(_8798_), .C(_8797_), .Y(_8799_) );
NAND2X1 NAND2X1_1648 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf1_), .B(_12588_), .Y(_8800_) );
OR2X2 OR2X2_288 ( .gnd(gnd), .vdd(vdd), .A(_12588_), .B(bloque_datos_24_bF_buf0_), .Y(_8801_) );
NAND2X1 NAND2X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .B(_8801_), .Y(_8802_) );
INVX2 INVX2_435 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .Y(_8803_) );
XNOR2X1 XNOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_10697_), .B(_8803_), .Y(_8804_) );
NAND3X1 NAND3X1_2851 ( .gnd(gnd), .vdd(vdd), .A(_8804_), .B(_8795_), .C(_8799_), .Y(_8805_) );
AOI21X1 AOI21X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_8798_), .B(_8797_), .C(_8796_), .Y(_8806_) );
AOI21X1 AOI21X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_8794_), .B(_8791_), .C(_12510_), .Y(_8807_) );
INVX1 INVX1_1750 ( .gnd(gnd), .vdd(vdd), .A(_8804_), .Y(_8808_) );
OAI21X1 OAI21X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_8806_), .B(_8807_), .C(_8808_), .Y(_8809_) );
AOI21X1 AOI21X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_8809_), .C(bloque_datos_52_bF_buf2_), .Y(_8810_) );
INVX1 INVX1_1751 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf1_), .Y(_8811_) );
NAND3X1 NAND3X1_2852 ( .gnd(gnd), .vdd(vdd), .A(_8808_), .B(_8795_), .C(_8799_), .Y(_8812_) );
OAI21X1 OAI21X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_8806_), .B(_8807_), .C(_8804_), .Y(_8813_) );
AOI21X1 AOI21X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_8813_), .C(_8811_), .Y(_8814_) );
OAI21X1 OAI21X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_8810_), .B(_8814_), .C(_12507_), .Y(_8815_) );
INVX2 INVX2_436 ( .gnd(gnd), .vdd(vdd), .A(_12507_), .Y(_8816_) );
NAND3X1 NAND3X1_2853 ( .gnd(gnd), .vdd(vdd), .A(_8811_), .B(_8812_), .C(_8813_), .Y(_8817_) );
NAND3X1 NAND3X1_2854 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf0_), .B(_8805_), .C(_8809_), .Y(_8818_) );
NAND3X1 NAND3X1_2855 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8817_), .C(_8818_), .Y(_8819_) );
NAND3X1 NAND3X1_2856 ( .gnd(gnd), .vdd(vdd), .A(_8819_), .B(_12505_), .C(_8815_), .Y(_8820_) );
OAI21X1 OAI21X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_12346_), .B(_12342_), .C(_12337_), .Y(_8821_) );
OAI21X1 OAI21X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_8810_), .B(_8814_), .C(_8816_), .Y(_8822_) );
NAND3X1 NAND3X1_2857 ( .gnd(gnd), .vdd(vdd), .A(_12507_), .B(_8817_), .C(_8818_), .Y(_8823_) );
NAND3X1 NAND3X1_2858 ( .gnd(gnd), .vdd(vdd), .A(_8823_), .B(_8822_), .C(_8821_), .Y(_8824_) );
NAND2X1 NAND2X1_1650 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf1_), .B(_8802_), .Y(_8825_) );
OR2X2 OR2X2_289 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(bloque_datos_40_bF_buf0_), .Y(_8826_) );
NAND2X1 NAND2X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_8826_), .Y(_8827_) );
INVX2 INVX2_437 ( .gnd(gnd), .vdd(vdd), .A(_8827_), .Y(_8828_) );
XNOR2X1 XNOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_10730_), .B(_8828_), .Y(_8829_) );
NAND3X1 NAND3X1_2859 ( .gnd(gnd), .vdd(vdd), .A(_8829_), .B(_8820_), .C(_8824_), .Y(_8830_) );
AOI21X1 AOI21X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_8823_), .B(_8822_), .C(_8821_), .Y(_8831_) );
AOI21X1 AOI21X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_8819_), .B(_8815_), .C(_12505_), .Y(_8832_) );
INVX1 INVX1_1752 ( .gnd(gnd), .vdd(vdd), .A(_8829_), .Y(_8833_) );
OAI21X1 OAI21X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_8831_), .B(_8832_), .C(_8833_), .Y(_8834_) );
AOI21X1 AOI21X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_8830_), .B(_8834_), .C(bloque_datos_68_bF_buf1_), .Y(_8835_) );
INVX1 INVX1_1753 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf0_), .Y(_8836_) );
NAND3X1 NAND3X1_2860 ( .gnd(gnd), .vdd(vdd), .A(_8833_), .B(_8820_), .C(_8824_), .Y(_8837_) );
OAI21X1 OAI21X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_8831_), .B(_8832_), .C(_8829_), .Y(_8838_) );
AOI21X1 AOI21X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_8837_), .B(_8838_), .C(_8836_), .Y(_8839_) );
OAI21X1 OAI21X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_8835_), .B(_8839_), .C(_12504_), .Y(_8840_) );
NAND3X1 NAND3X1_2861 ( .gnd(gnd), .vdd(vdd), .A(_8836_), .B(_8837_), .C(_8838_), .Y(_8841_) );
NAND3X1 NAND3X1_2862 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf3_), .B(_8830_), .C(_8834_), .Y(_8842_) );
NAND3X1 NAND3X1_2863 ( .gnd(gnd), .vdd(vdd), .A(_12353_), .B(_8841_), .C(_8842_), .Y(_8843_) );
NAND3X1 NAND3X1_2864 ( .gnd(gnd), .vdd(vdd), .A(_12503_), .B(_8843_), .C(_8840_), .Y(_8844_) );
INVX1 INVX1_1754 ( .gnd(gnd), .vdd(vdd), .A(_12271_), .Y(_8845_) );
AOI21X1 AOI21X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_12348_), .B(_12351_), .C(_12140_), .Y(_8846_) );
OAI21X1 OAI21X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_8846_), .B(_8845_), .C(_12352_), .Y(_8847_) );
OAI21X1 OAI21X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_8835_), .B(_8839_), .C(_12353_), .Y(_8848_) );
NAND3X1 NAND3X1_2865 ( .gnd(gnd), .vdd(vdd), .A(_12504_), .B(_8841_), .C(_8842_), .Y(_8849_) );
NAND3X1 NAND3X1_2866 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .B(_8849_), .C(_8848_), .Y(_8850_) );
NAND2X1 NAND2X1_1652 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf1_), .B(_8827_), .Y(_8851_) );
OR2X2 OR2X2_290 ( .gnd(gnd), .vdd(vdd), .A(_8827_), .B(bloque_datos_56_bF_buf0_), .Y(_8852_) );
NAND2X1 NAND2X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_8851_), .B(_8852_), .Y(_8853_) );
INVX2 INVX2_438 ( .gnd(gnd), .vdd(vdd), .A(_8853_), .Y(_8854_) );
XNOR2X1 XNOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_10763_), .B(_8854_), .Y(_8855_) );
NAND3X1 NAND3X1_2867 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_8844_), .C(_8850_), .Y(_8856_) );
AOI21X1 AOI21X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_8849_), .B(_8848_), .C(_8847_), .Y(_8857_) );
AOI21X1 AOI21X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_8843_), .B(_8840_), .C(_12503_), .Y(_8858_) );
INVX1 INVX1_1755 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .Y(_8859_) );
OAI21X1 OAI21X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_8858_), .C(_8859_), .Y(_8860_) );
AOI21X1 AOI21X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_8856_), .B(_8860_), .C(bloque_datos_84_bF_buf2_), .Y(_8861_) );
INVX1 INVX1_1756 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf1_), .Y(_8862_) );
NAND3X1 NAND3X1_2868 ( .gnd(gnd), .vdd(vdd), .A(_8859_), .B(_8844_), .C(_8850_), .Y(_8863_) );
OAI21X1 OAI21X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_8858_), .C(_8855_), .Y(_8864_) );
AOI21X1 AOI21X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_8863_), .B(_8864_), .C(_8862_), .Y(_8865_) );
OAI21X1 OAI21X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .B(_8865_), .C(_12501_), .Y(_8866_) );
NAND3X1 NAND3X1_2869 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .B(_8863_), .C(_8864_), .Y(_8867_) );
NAND3X1 NAND3X1_2870 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf0_), .B(_8856_), .C(_8860_), .Y(_8868_) );
NAND3X1 NAND3X1_2871 ( .gnd(gnd), .vdd(vdd), .A(_12365_), .B(_8867_), .C(_8868_), .Y(_8869_) );
NAND3X1 NAND3X1_2872 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_8869_), .C(_12500_), .Y(_8870_) );
NAND2X1 NAND2X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_12363_), .B(_12369_), .Y(_8871_) );
OAI21X1 OAI21X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .B(_8865_), .C(_12365_), .Y(_8872_) );
NAND3X1 NAND3X1_2873 ( .gnd(gnd), .vdd(vdd), .A(_12501_), .B(_8867_), .C(_8868_), .Y(_8873_) );
NAND3X1 NAND3X1_2874 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8873_), .C(_8872_), .Y(_8874_) );
NOR2X1 NOR2X1_963 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf2_), .B(_8854_), .Y(_8875_) );
NAND2X1 NAND2X1_1655 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf1_), .B(_8854_), .Y(_8876_) );
INVX1 INVX1_1757 ( .gnd(gnd), .vdd(vdd), .A(_8876_), .Y(_8877_) );
NOR2X1 NOR2X1_964 ( .gnd(gnd), .vdd(vdd), .A(_8875_), .B(_8877_), .Y(_8878_) );
XOR2X1 XOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_10796_), .B(_8878_), .Y(_8879_) );
NAND3X1 NAND3X1_2875 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(_8874_), .C(_8870_), .Y(_8880_) );
AOI21X1 AOI21X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_8873_), .B(_8872_), .C(_8871_), .Y(_8881_) );
AOI21X1 AOI21X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_8869_), .B(_8866_), .C(_12500_), .Y(_8882_) );
INVX1 INVX1_1758 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .Y(_8883_) );
OAI21X1 OAI21X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_8881_), .B(_8882_), .C(_8883_), .Y(_8884_) );
AOI21X1 AOI21X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_8884_), .C(module_2_W_132_), .Y(_8885_) );
INVX1 INVX1_1759 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_132_), .Y(_8886_) );
NAND3X1 NAND3X1_2876 ( .gnd(gnd), .vdd(vdd), .A(_8883_), .B(_8874_), .C(_8870_), .Y(_8887_) );
OAI21X1 OAI21X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_8881_), .B(_8882_), .C(_8879_), .Y(_8888_) );
AOI21X1 AOI21X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_8887_), .B(_8888_), .C(_8886_), .Y(_8889_) );
OAI21X1 OAI21X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_8885_), .B(_8889_), .C(_12371_), .Y(_8890_) );
INVX2 INVX2_439 ( .gnd(gnd), .vdd(vdd), .A(_12371_), .Y(_8891_) );
NAND3X1 NAND3X1_2877 ( .gnd(gnd), .vdd(vdd), .A(_8886_), .B(_8887_), .C(_8888_), .Y(_8892_) );
NAND3X1 NAND3X1_2878 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_132_), .B(_8880_), .C(_8884_), .Y(_8893_) );
NAND3X1 NAND3X1_2879 ( .gnd(gnd), .vdd(vdd), .A(_8891_), .B(_8892_), .C(_8893_), .Y(_8894_) );
AOI21X1 AOI21X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_8894_), .B(_8890_), .C(_12499_), .Y(_8895_) );
AND2X2 AND2X2_278 ( .gnd(gnd), .vdd(vdd), .A(_12378_), .B(_12375_), .Y(_8896_) );
OAI21X1 OAI21X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_8885_), .B(_8889_), .C(_8891_), .Y(_8897_) );
NAND3X1 NAND3X1_2880 ( .gnd(gnd), .vdd(vdd), .A(_12371_), .B(_8892_), .C(_8893_), .Y(_8898_) );
AOI21X1 AOI21X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_8898_), .B(_8897_), .C(_8896_), .Y(_8899_) );
NAND2X1 NAND2X1_1656 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf4_), .B(_8878_), .Y(_8900_) );
OR2X2 OR2X2_291 ( .gnd(gnd), .vdd(vdd), .A(_8878_), .B(bloque_datos_88_bF_buf3_), .Y(_8901_) );
NAND2X1 NAND2X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_8900_), .B(_8901_), .Y(_8902_) );
OAI21X1 OAI21X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_8895_), .B(_8899_), .C(_8902_), .Y(_8903_) );
AOI21X1 AOI21X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_8892_), .B(_8893_), .C(_8891_), .Y(_8904_) );
NOR3X1 NOR3X1_370 ( .gnd(gnd), .vdd(vdd), .A(_8885_), .B(_12371_), .C(_8889_), .Y(_8905_) );
OAI21X1 OAI21X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_8905_), .B(_8904_), .C(_8896_), .Y(_8906_) );
NAND3X1 NAND3X1_2881 ( .gnd(gnd), .vdd(vdd), .A(_12499_), .B(_8894_), .C(_8890_), .Y(_8907_) );
INVX2 INVX2_440 ( .gnd(gnd), .vdd(vdd), .A(_8902_), .Y(_8908_) );
NAND3X1 NAND3X1_2882 ( .gnd(gnd), .vdd(vdd), .A(_8907_), .B(_8908_), .C(_8906_), .Y(_8909_) );
NAND2X1 NAND2X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_8909_), .Y(_8910_) );
NAND3X1 NAND3X1_2883 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_148_), .B(_10829_), .C(_8910_), .Y(_8911_) );
INVX1 INVX1_1760 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_148_), .Y(_8912_) );
AOI21X1 AOI21X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_8907_), .B(_8906_), .C(_8902_), .Y(_8913_) );
NAND2X1 NAND2X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_8907_), .B(_8906_), .Y(_8914_) );
OAI21X1 OAI21X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_8914_), .B(_8908_), .C(_10829_), .Y(_8915_) );
OAI21X1 OAI21X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_8915_), .B(_8913_), .C(_8912_), .Y(_8916_) );
AOI21X1 AOI21X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_8916_), .C(_12384_), .Y(_8917_) );
OAI21X1 OAI21X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_8915_), .B(_8913_), .C(module_2_W_148_), .Y(_8918_) );
NAND3X1 NAND3X1_2884 ( .gnd(gnd), .vdd(vdd), .A(_8912_), .B(_10829_), .C(_8910_), .Y(_8919_) );
AOI21X1 AOI21X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_8919_), .B(_8918_), .C(_12383_), .Y(_8920_) );
OAI21X1 OAI21X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_8920_), .B(_8917_), .C(_12498_), .Y(_8921_) );
NAND2X1 NAND2X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_12385_), .B(_12389_), .Y(_8922_) );
NAND3X1 NAND3X1_2885 ( .gnd(gnd), .vdd(vdd), .A(_12383_), .B(_8919_), .C(_8918_), .Y(_8923_) );
NAND3X1 NAND3X1_2886 ( .gnd(gnd), .vdd(vdd), .A(_12384_), .B(_8911_), .C(_8916_), .Y(_8924_) );
NAND3X1 NAND3X1_2887 ( .gnd(gnd), .vdd(vdd), .A(_8922_), .B(_8923_), .C(_8924_), .Y(_8925_) );
NAND2X1 NAND2X1_1661 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_136_), .B(_8902_), .Y(_8926_) );
OR2X2 OR2X2_292 ( .gnd(gnd), .vdd(vdd), .A(_8902_), .B(module_2_W_136_), .Y(_8927_) );
NAND2X1 NAND2X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_8926_), .B(_8927_), .Y(_8928_) );
NAND3X1 NAND3X1_2888 ( .gnd(gnd), .vdd(vdd), .A(_8925_), .B(_8928_), .C(_8921_), .Y(_8929_) );
NAND2X1 NAND2X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_8925_), .B(_8921_), .Y(_8930_) );
INVX2 INVX2_441 ( .gnd(gnd), .vdd(vdd), .A(_8928_), .Y(_8931_) );
AOI21X1 AOI21X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_8931_), .B(_8930_), .C(_11114_), .Y(_8932_) );
NAND3X1 NAND3X1_2889 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_164_), .B(_8929_), .C(_8932_), .Y(_8933_) );
INVX1 INVX1_1761 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_164_), .Y(_8934_) );
AOI21X1 AOI21X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .B(_8924_), .C(_8922_), .Y(_8935_) );
NAND3X1 NAND3X1_2890 ( .gnd(gnd), .vdd(vdd), .A(_12383_), .B(_8911_), .C(_8916_), .Y(_8936_) );
NAND3X1 NAND3X1_2891 ( .gnd(gnd), .vdd(vdd), .A(_12384_), .B(_8919_), .C(_8918_), .Y(_8937_) );
AOI21X1 AOI21X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_8936_), .B(_8937_), .C(_12498_), .Y(_8938_) );
OAI21X1 OAI21X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_8935_), .B(_8938_), .C(_8931_), .Y(_8939_) );
NAND3X1 NAND3X1_2892 ( .gnd(gnd), .vdd(vdd), .A(_10862_), .B(_8929_), .C(_8939_), .Y(_8940_) );
NAND2X1 NAND2X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_8934_), .B(_8940_), .Y(_8941_) );
AOI21X1 AOI21X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_8941_), .B(_8933_), .C(_12394_), .Y(_8942_) );
INVX1 INVX1_1762 ( .gnd(gnd), .vdd(vdd), .A(_12394_), .Y(_8943_) );
NAND2X1 NAND2X1_1665 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_164_), .B(_8940_), .Y(_8944_) );
NAND3X1 NAND3X1_2893 ( .gnd(gnd), .vdd(vdd), .A(_8934_), .B(_8929_), .C(_8932_), .Y(_8945_) );
AOI21X1 AOI21X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_8945_), .C(_8943_), .Y(_8946_) );
OAI21X1 OAI21X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_8946_), .B(_8942_), .C(_12497_), .Y(_8947_) );
NAND3X1 NAND3X1_2894 ( .gnd(gnd), .vdd(vdd), .A(_8943_), .B(_8944_), .C(_8945_), .Y(_8948_) );
NAND3X1 NAND3X1_2895 ( .gnd(gnd), .vdd(vdd), .A(_12394_), .B(_8941_), .C(_8933_), .Y(_8949_) );
NAND3X1 NAND3X1_2896 ( .gnd(gnd), .vdd(vdd), .A(_12496_), .B(_8948_), .C(_8949_), .Y(_8950_) );
NAND2X1 NAND2X1_1666 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_152_), .B(_8928_), .Y(_8951_) );
OR2X2 OR2X2_293 ( .gnd(gnd), .vdd(vdd), .A(_8928_), .B(module_2_W_152_), .Y(_8952_) );
NAND2X1 NAND2X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_8951_), .B(_8952_), .Y(_8953_) );
NAND3X1 NAND3X1_2897 ( .gnd(gnd), .vdd(vdd), .A(_8950_), .B(_8953_), .C(_8947_), .Y(_8954_) );
AOI21X1 AOI21X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_8950_), .B(_8947_), .C(_8953_), .Y(_8955_) );
NOR2X1 NOR2X1_965 ( .gnd(gnd), .vdd(vdd), .A(_11092_), .B(_8955_), .Y(_8956_) );
NAND3X1 NAND3X1_2898 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_180_), .B(_8954_), .C(_8956_), .Y(_8957_) );
INVX1 INVX1_1763 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_180_), .Y(_8958_) );
NAND2X1 NAND2X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_10895_), .B(_8954_), .Y(_8959_) );
OAI21X1 OAI21X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_8959_), .B(_8955_), .C(_8958_), .Y(_8960_) );
AOI21X1 AOI21X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_8960_), .B(_8957_), .C(_12407_), .Y(_8961_) );
OAI21X1 OAI21X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_8959_), .B(_8955_), .C(module_2_W_180_), .Y(_8962_) );
NAND3X1 NAND3X1_2899 ( .gnd(gnd), .vdd(vdd), .A(_8958_), .B(_8954_), .C(_8956_), .Y(_8963_) );
AOI21X1 AOI21X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_8962_), .B(_8963_), .C(_12406_), .Y(_8964_) );
OAI21X1 OAI21X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_8964_), .B(_8961_), .C(_12494_), .Y(_8965_) );
OAI21X1 OAI21X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_12414_), .B(_12261_), .C(_12408_), .Y(_8966_) );
NAND3X1 NAND3X1_2900 ( .gnd(gnd), .vdd(vdd), .A(_12406_), .B(_8962_), .C(_8963_), .Y(_8967_) );
NAND3X1 NAND3X1_2901 ( .gnd(gnd), .vdd(vdd), .A(_12407_), .B(_8960_), .C(_8957_), .Y(_8968_) );
NAND3X1 NAND3X1_2902 ( .gnd(gnd), .vdd(vdd), .A(_8967_), .B(_8966_), .C(_8968_), .Y(_8969_) );
NAND2X1 NAND2X1_1669 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_168_), .B(_8953_), .Y(_8970_) );
OR2X2 OR2X2_294 ( .gnd(gnd), .vdd(vdd), .A(_8953_), .B(module_2_W_168_), .Y(_8971_) );
NAND2X1 NAND2X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_8970_), .B(_8971_), .Y(_8972_) );
NAND3X1 NAND3X1_2903 ( .gnd(gnd), .vdd(vdd), .A(_8969_), .B(_8972_), .C(_8965_), .Y(_8973_) );
NAND2X1 NAND2X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_8969_), .B(_8965_), .Y(_8974_) );
INVX2 INVX2_442 ( .gnd(gnd), .vdd(vdd), .A(_8972_), .Y(_8975_) );
AOI21X1 AOI21X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_8975_), .B(_8974_), .C(_11059_), .Y(_8976_) );
NAND3X1 NAND3X1_2904 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_196_), .B(_8973_), .C(_8976_), .Y(_8977_) );
INVX1 INVX1_1764 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_196_), .Y(_8978_) );
AOI21X1 AOI21X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_8967_), .B(_8968_), .C(_8966_), .Y(_8979_) );
NOR3X1 NOR3X1_371 ( .gnd(gnd), .vdd(vdd), .A(_8961_), .B(_12494_), .C(_8964_), .Y(_8980_) );
OAI21X1 OAI21X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_8980_), .B(_8979_), .C(_8975_), .Y(_8981_) );
NAND3X1 NAND3X1_2905 ( .gnd(gnd), .vdd(vdd), .A(_10928_), .B(_8973_), .C(_8981_), .Y(_8982_) );
NAND2X1 NAND2X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_8978_), .B(_8982_), .Y(_8983_) );
AOI21X1 AOI21X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_8977_), .B(_8983_), .C(_12419_), .Y(_8984_) );
INVX1 INVX1_1765 ( .gnd(gnd), .vdd(vdd), .A(_12412_), .Y(_8985_) );
NAND2X1 NAND2X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_12415_), .B(_8985_), .Y(_8986_) );
NOR2X1 NOR2X1_966 ( .gnd(gnd), .vdd(vdd), .A(_12260_), .B(_8986_), .Y(_8987_) );
NAND2X1 NAND2X1_1674 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_196_), .B(_8982_), .Y(_8988_) );
NAND3X1 NAND3X1_2906 ( .gnd(gnd), .vdd(vdd), .A(_8978_), .B(_8973_), .C(_8976_), .Y(_8989_) );
AOI21X1 AOI21X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_8989_), .B(_8988_), .C(_8987_), .Y(_8990_) );
OAI21X1 OAI21X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_8984_), .B(_8990_), .C(_12492_), .Y(_8991_) );
OAI21X1 OAI21X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_12422_), .B(_12258_), .C(_12421_), .Y(_8992_) );
NAND3X1 NAND3X1_2907 ( .gnd(gnd), .vdd(vdd), .A(_8987_), .B(_8989_), .C(_8988_), .Y(_8993_) );
NAND3X1 NAND3X1_2908 ( .gnd(gnd), .vdd(vdd), .A(_12419_), .B(_8977_), .C(_8983_), .Y(_8994_) );
NAND3X1 NAND3X1_2909 ( .gnd(gnd), .vdd(vdd), .A(_8993_), .B(_8994_), .C(_8992_), .Y(_8995_) );
NAND2X1 NAND2X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_8995_), .B(_8991_), .Y(_8996_) );
NAND2X1 NAND2X1_1676 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_184_), .B(_8972_), .Y(_8997_) );
OR2X2 OR2X2_295 ( .gnd(gnd), .vdd(vdd), .A(_8972_), .B(module_2_W_184_), .Y(_8998_) );
NAND2X1 NAND2X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_8997_), .B(_8998_), .Y(_8999_) );
INVX2 INVX2_443 ( .gnd(gnd), .vdd(vdd), .A(_8999_), .Y(_9000_) );
OR2X2 OR2X2_296 ( .gnd(gnd), .vdd(vdd), .A(_8996_), .B(_9000_), .Y(_9001_) );
AOI21X1 AOI21X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_8995_), .B(_8991_), .C(_8999_), .Y(_9002_) );
NOR2X1 NOR2X1_967 ( .gnd(gnd), .vdd(vdd), .A(_11038_), .B(_9002_), .Y(_9003_) );
NAND3X1 NAND3X1_2910 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_212_), .B(_9001_), .C(_9003_), .Y(_9004_) );
INVX1 INVX1_1766 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_212_), .Y(_9005_) );
OAI21X1 OAI21X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_8996_), .B(_9000_), .C(_10961_), .Y(_9006_) );
OAI21X1 OAI21X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_9006_), .B(_9002_), .C(_9005_), .Y(_9007_) );
AOI21X1 AOI21X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_9007_), .B(_9004_), .C(_12437_), .Y(_9008_) );
OAI21X1 OAI21X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_9006_), .B(_9002_), .C(module_2_W_212_), .Y(_9009_) );
NAND3X1 NAND3X1_2911 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(_9001_), .C(_9003_), .Y(_9010_) );
AOI21X1 AOI21X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_9009_), .B(_9010_), .C(_12434_), .Y(_9011_) );
OAI21X1 OAI21X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_9008_), .B(_9011_), .C(_12490_), .Y(_9012_) );
NAND3X1 NAND3X1_2912 ( .gnd(gnd), .vdd(vdd), .A(_12215_), .B(_12429_), .C(_12437_), .Y(_9013_) );
OAI21X1 OAI21X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_12441_), .B(_12438_), .C(_9013_), .Y(_9014_) );
NAND3X1 NAND3X1_2913 ( .gnd(gnd), .vdd(vdd), .A(_12434_), .B(_9009_), .C(_9010_), .Y(_9015_) );
NAND3X1 NAND3X1_2914 ( .gnd(gnd), .vdd(vdd), .A(_12437_), .B(_9007_), .C(_9004_), .Y(_9016_) );
INVX1 INVX1_1767 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_0_), .Y(_12772_) );
INVX4 INVX4_11 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf0), .Y(_12773_) );
NAND2X1 NAND2X1_1678 ( .gnd(gnd), .vdd(vdd), .A(nonce_iniciales[64]), .B(_12773_), .Y(_12593_) );
OAI21X1 OAI21X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_12772_), .B(_12773_), .C(_12593_), .Y(_12592__0_) );
INVX1 INVX1_1768 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_1_), .Y(_12594_) );
NAND2X1 NAND2X1_1679 ( .gnd(gnd), .vdd(vdd), .A(nonce_iniciales[65]), .B(_12773_), .Y(_12595_) );
OAI21X1 OAI21X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_12773_), .B(_12594_), .C(_12595_), .Y(_12592__1_) );
NAND2X1 NAND2X1_1680 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_5_), .B(module_2_W_4_), .Y(_12596_) );
NAND2X1 NAND2X1_1681 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_7_), .B(module_2_W_6_), .Y(_12597_) );
NOR2X1 NOR2X1_968 ( .gnd(gnd), .vdd(vdd), .A(_12596_), .B(_12597_), .Y(_12598_) );
NAND2X1 NAND2X1_1682 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_25_), .B(module_2_W_24_), .Y(_12599_) );
NAND2X1 NAND2X1_1683 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_27_), .B(module_2_W_26_), .Y(_12600_) );
NOR2X1 NOR2X1_969 ( .gnd(gnd), .vdd(vdd), .A(_12599_), .B(_12600_), .Y(_12601_) );
INVX1 INVX1_1769 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_2_), .Y(_12602_) );
OAI21X1 OAI21X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_12772_), .B(_12594_), .C(_12602_), .Y(_12603_) );
NAND3X1 NAND3X1_2915 ( .gnd(gnd), .vdd(vdd), .A(_12603_), .B(_12598_), .C(_12601_), .Y(_12604_) );
INVX1 INVX1_1770 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_29_), .Y(_12605_) );
INVX1 INVX1_1771 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_28_), .Y(_12606_) );
NOR2X1 NOR2X1_970 ( .gnd(gnd), .vdd(vdd), .A(_12605_), .B(_12606_), .Y(_12607_) );
INVX1 INVX1_1772 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_31_), .Y(_12608_) );
INVX1 INVX1_1773 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_30_), .Y(_12609_) );
NOR2X1 NOR2X1_971 ( .gnd(gnd), .vdd(vdd), .A(_12608_), .B(_12609_), .Y(_12610_) );
NAND3X1 NAND3X1_2916 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_3_), .B(_12607_), .C(_12610_), .Y(_12611_) );
NOR2X1 NOR2X1_972 ( .gnd(gnd), .vdd(vdd), .A(_12611_), .B(_12604_), .Y(_12612_) );
NAND2X1 NAND2X1_1684 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_17_), .B(module_2_W_16_), .Y(_12613_) );
NAND2X1 NAND2X1_1685 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_19_), .B(module_2_W_18_), .Y(_12614_) );
NOR2X1 NOR2X1_973 ( .gnd(gnd), .vdd(vdd), .A(_12613_), .B(_12614_), .Y(_12615_) );
NAND2X1 NAND2X1_1686 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_22_), .B(module_2_W_21_), .Y(_12616_) );
NAND2X1 NAND2X1_1687 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_23_), .B(module_2_W_20_), .Y(_12617_) );
NOR2X1 NOR2X1_974 ( .gnd(gnd), .vdd(vdd), .A(_12616_), .B(_12617_), .Y(_12618_) );
NAND2X1 NAND2X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_12615_), .B(_12618_), .Y(_12619_) );
NAND2X1 NAND2X1_1689 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_9_), .B(module_2_W_8_), .Y(_12620_) );
NAND2X1 NAND2X1_1690 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_11_), .B(module_2_W_10_), .Y(_12621_) );
NOR2X1 NOR2X1_975 ( .gnd(gnd), .vdd(vdd), .A(_12620_), .B(_12621_), .Y(_12622_) );
NAND2X1 NAND2X1_1691 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_15_), .B(module_2_W_14_), .Y(_12623_) );
NAND2X1 NAND2X1_1692 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_13_), .B(module_2_W_12_), .Y(_12624_) );
NOR2X1 NOR2X1_976 ( .gnd(gnd), .vdd(vdd), .A(_12623_), .B(_12624_), .Y(_12625_) );
NAND2X1 NAND2X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_12622_), .B(_12625_), .Y(_12626_) );
NOR2X1 NOR2X1_977 ( .gnd(gnd), .vdd(vdd), .A(_12619_), .B(_12626_), .Y(_12627_) );
AOI21X1 AOI21X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_12627_), .B(_12612_), .C(_12773_), .Y(_12628_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_2_), .B(nonce_iniciales[66]), .S(inicio_bF_buf0), .Y(_12629_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_2_), .B(_12629_), .S(_12628__bF_buf1), .Y(_12592__2_) );
NAND2X1 NAND2X1_1694 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_2_), .B(module_2_W_3_), .Y(_12630_) );
INVX1 INVX1_1774 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_3_), .Y(_12631_) );
NAND2X1 NAND2X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_12602_), .B(_12631_), .Y(_12632_) );
NAND2X1 NAND2X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_12630_), .B(_12632_), .Y(_12633_) );
NOR2X1 NOR2X1_978 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf0), .B(nonce_iniciales[67]), .Y(_12634_) );
AOI21X1 AOI21X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_12633_), .B(_12628__bF_buf0), .C(_12634_), .Y(_12592__3_) );
XOR2X1 XOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_12630_), .B(module_2_W_4_), .Y(_12635_) );
NOR2X1 NOR2X1_979 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf0), .B(nonce_iniciales[68]), .Y(_12636_) );
AOI21X1 AOI21X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_12635_), .B(_12628__bF_buf1), .C(_12636_), .Y(_12592__4_) );
AND2X2 AND2X2_279 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_2_), .B(module_2_W_3_), .Y(_12637_) );
NAND2X1 NAND2X1_1697 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_4_), .B(_12637_), .Y(_12638_) );
XOR2X1 XOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_12638_), .B(module_2_W_5_), .Y(_12639_) );
NOR2X1 NOR2X1_980 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[69]), .Y(_12640_) );
AOI21X1 AOI21X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_12639_), .B(_12628__bF_buf0), .C(_12640_), .Y(_12592__5_) );
NOR2X1 NOR2X1_981 ( .gnd(gnd), .vdd(vdd), .A(_12596_), .B(_12630_), .Y(_12641_) );
XNOR2X1 XNOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_12641_), .B(module_2_W_6_), .Y(_12642_) );
NOR2X1 NOR2X1_982 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[70]), .Y(_12643_) );
AOI21X1 AOI21X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_12642_), .B(_12628__bF_buf1), .C(_12643_), .Y(_12592__6_) );
NOR2X1 NOR2X1_983 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[71]), .Y(_12644_) );
NAND2X1 NAND2X1_1698 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_6_), .B(_12641_), .Y(_12645_) );
XOR2X1 XOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_12645_), .B(module_2_W_7_), .Y(_12646_) );
AOI21X1 AOI21X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_12646_), .B(_12628__bF_buf1), .C(_12644_), .Y(_12592__7_) );
NOR3X1 NOR3X1_372 ( .gnd(gnd), .vdd(vdd), .A(_12596_), .B(_12597_), .C(_12630_), .Y(_12647_) );
XNOR2X1 XNOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_12647_), .B(module_2_W_8_), .Y(_12648_) );
NOR2X1 NOR2X1_984 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[72]), .Y(_12649_) );
AOI21X1 AOI21X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_12648_), .B(_12628__bF_buf2), .C(_12649_), .Y(_12592__8_) );
AND2X2 AND2X2_280 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_5_), .B(module_2_W_4_), .Y(_12650_) );
AND2X2 AND2X2_281 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_7_), .B(module_2_W_6_), .Y(_12651_) );
NAND3X1 NAND3X1_2917 ( .gnd(gnd), .vdd(vdd), .A(_12650_), .B(_12651_), .C(_12637_), .Y(_12652_) );
INVX1 INVX1_1775 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_9_), .Y(_12653_) );
INVX1 INVX1_1776 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_8_), .Y(_12654_) );
OAI21X1 OAI21X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_12652_), .B(_12654_), .C(_12653_), .Y(_12655_) );
OAI21X1 OAI21X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_12620_), .B(_12652_), .C(_12655_), .Y(_12656_) );
NOR2X1 NOR2X1_985 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[73]), .Y(_12657_) );
AOI21X1 AOI21X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_12656_), .B(_12628__bF_buf2), .C(_12657_), .Y(_12592__9_) );
NOR2X1 NOR2X1_986 ( .gnd(gnd), .vdd(vdd), .A(_12620_), .B(_12652_), .Y(_12658_) );
XNOR2X1 XNOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_12658_), .B(module_2_W_10_), .Y(_12659_) );
NOR2X1 NOR2X1_987 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[74]), .Y(_12660_) );
AOI21X1 AOI21X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_12659_), .B(_12628__bF_buf1), .C(_12660_), .Y(_12592__10_) );
NOR2X1 NOR2X1_988 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[75]), .Y(_12661_) );
NAND2X1 NAND2X1_1699 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_10_), .B(_12658_), .Y(_12662_) );
OR2X2 OR2X2_297 ( .gnd(gnd), .vdd(vdd), .A(_12662_), .B(module_2_W_11_), .Y(_12663_) );
NAND2X1 NAND2X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_12627_), .B(_12612_), .Y(_12664_) );
NAND2X1 NAND2X1_1701 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf0), .B(_12664_), .Y(_12665_) );
AOI21X1 AOI21X1_1795 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_11_), .B(_12662_), .C(_12665_), .Y(_12666_) );
AOI21X1 AOI21X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_12663_), .B(_12666_), .C(_12661_), .Y(_12592__11_) );
INVX2 INVX2_444 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_12_), .Y(_12667_) );
NAND2X1 NAND2X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_12622_), .B(_12647_), .Y(_12668_) );
XNOR2X1 XNOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_12668_), .B(_12667_), .Y(_12669_) );
NOR2X1 NOR2X1_989 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[76]), .Y(_12670_) );
AOI21X1 AOI21X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_12669_), .B(_12628__bF_buf2), .C(_12670_), .Y(_12592__12_) );
NOR2X1 NOR2X1_990 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[77]), .Y(_12671_) );
INVX1 INVX1_1777 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_13_), .Y(_12672_) );
NAND3X1 NAND3X1_2918 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_11_), .B(module_2_W_10_), .C(_12658_), .Y(_12673_) );
NOR2X1 NOR2X1_991 ( .gnd(gnd), .vdd(vdd), .A(_12667_), .B(_12673_), .Y(_12674_) );
NAND2X1 NAND2X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_12672_), .B(_12674_), .Y(_12675_) );
OAI21X1 OAI21X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_12668_), .B(_12667_), .C(module_2_W_13_), .Y(_12676_) );
AND2X2 AND2X2_282 ( .gnd(gnd), .vdd(vdd), .A(_12628__bF_buf2), .B(_12676_), .Y(_12677_) );
AOI21X1 AOI21X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_12675_), .B(_12677_), .C(_12671_), .Y(_12592__13_) );
INVX2 INVX2_445 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_14_), .Y(_12678_) );
OR2X2 OR2X2_298 ( .gnd(gnd), .vdd(vdd), .A(_12668_), .B(_12624_), .Y(_12679_) );
XNOR2X1 XNOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_12679_), .B(_12678_), .Y(_12680_) );
NOR2X1 NOR2X1_992 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[78]), .Y(_12681_) );
AOI21X1 AOI21X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_12628__bF_buf2), .B(_12680_), .C(_12681_), .Y(_12592__14_) );
NOR2X1 NOR2X1_993 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[79]), .Y(_12682_) );
INVX1 INVX1_1778 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_15_), .Y(_12683_) );
NOR2X1 NOR2X1_994 ( .gnd(gnd), .vdd(vdd), .A(_12624_), .B(_12673_), .Y(_12684_) );
NAND3X1 NAND3X1_2919 ( .gnd(gnd), .vdd(vdd), .A(_12683_), .B(module_2_W_14_), .C(_12684_), .Y(_12685_) );
OAI21X1 OAI21X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_12679_), .B(_12678_), .C(module_2_W_15_), .Y(_12686_) );
AND2X2 AND2X2_283 ( .gnd(gnd), .vdd(vdd), .A(_12686_), .B(_12628__bF_buf2), .Y(_12687_) );
AOI21X1 AOI21X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_12685_), .B(_12687_), .C(_12682_), .Y(_12592__15_) );
OR2X2 OR2X2_299 ( .gnd(gnd), .vdd(vdd), .A(_12620_), .B(_12621_), .Y(_12688_) );
OR2X2 OR2X2_300 ( .gnd(gnd), .vdd(vdd), .A(_12623_), .B(_12624_), .Y(_12689_) );
NOR3X1 NOR3X1_373 ( .gnd(gnd), .vdd(vdd), .A(_12689_), .B(_12688_), .C(_12652_), .Y(_12690_) );
NAND2X1 NAND2X1_1704 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_16_), .B(_12690_), .Y(_12691_) );
INVX1 INVX1_1779 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_16_), .Y(_12692_) );
OAI21X1 OAI21X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_12626_), .B(_12652_), .C(_12692_), .Y(_12693_) );
NAND2X1 NAND2X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_12693_), .B(_12691_), .Y(_12694_) );
NOR2X1 NOR2X1_995 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf0), .B(nonce_iniciales[80]), .Y(_12695_) );
AOI21X1 AOI21X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_12628__bF_buf0), .B(_12694_), .C(_12695_), .Y(_12592__16_) );
NAND3X1 NAND3X1_2920 ( .gnd(gnd), .vdd(vdd), .A(_12622_), .B(_12625_), .C(_12647_), .Y(_12696_) );
NOR2X1 NOR2X1_996 ( .gnd(gnd), .vdd(vdd), .A(_12692_), .B(_12696_), .Y(_12697_) );
XNOR2X1 XNOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_12697_), .B(module_2_W_17_), .Y(_12698_) );
NOR2X1 NOR2X1_997 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf1), .B(nonce_iniciales[81]), .Y(_12699_) );
AOI21X1 AOI21X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_12628__bF_buf3), .B(_12698_), .C(_12699_), .Y(_12592__17_) );
INVX1 INVX1_1780 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_18_), .Y(_12700_) );
INVX1 INVX1_1781 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_17_), .Y(_12701_) );
OAI21X1 OAI21X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_12691_), .B(_12701_), .C(_12700_), .Y(_12702_) );
NAND3X1 NAND3X1_2921 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_18_), .B(module_2_W_17_), .C(_12697_), .Y(_12703_) );
NAND2X1 NAND2X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_12703_), .B(_12702_), .Y(_12704_) );
NOR2X1 NOR2X1_998 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf1), .B(nonce_iniciales[82]), .Y(_12705_) );
AOI21X1 AOI21X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_12628__bF_buf3), .B(_12704_), .C(_12705_), .Y(_12592__18_) );
NOR2X1 NOR2X1_999 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf1), .B(nonce_iniciales[83]), .Y(_12706_) );
OR2X2 OR2X2_301 ( .gnd(gnd), .vdd(vdd), .A(_12703_), .B(module_2_W_19_), .Y(_12707_) );
AOI21X1 AOI21X1_1804 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_19_), .B(_12703_), .C(_12665_), .Y(_12708_) );
AOI21X1 AOI21X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_12707_), .B(_12708_), .C(_12706_), .Y(_12592__19_) );
INVX1 INVX1_1782 ( .gnd(gnd), .vdd(vdd), .A(_12615_), .Y(_12709_) );
NOR2X1 NOR2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_12709_), .B(_12696_), .Y(_12710_) );
NAND2X1 NAND2X1_1707 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_20_), .B(_12710_), .Y(_12711_) );
INVX2 INVX2_446 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_20_), .Y(_12712_) );
OAI21X1 OAI21X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_12696_), .B(_12709_), .C(_12712_), .Y(_12713_) );
NAND2X1 NAND2X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_12713_), .B(_12711_), .Y(_12714_) );
NOR2X1 NOR2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf1), .B(nonce_iniciales[84]), .Y(_12715_) );
AOI21X1 AOI21X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_12628__bF_buf3), .B(_12714_), .C(_12715_), .Y(_12592__20_) );
INVX1 INVX1_1783 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_21_), .Y(_12716_) );
INVX1 INVX1_1784 ( .gnd(gnd), .vdd(vdd), .A(_12664_), .Y(_12717_) );
NAND2X1 NAND2X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_12615_), .B(_12690_), .Y(_12718_) );
NOR2X1 NOR2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_12712_), .B(_12718_), .Y(_12719_) );
AOI21X1 AOI21X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_12716_), .B(_12719_), .C(_12717_), .Y(_12720_) );
AOI21X1 AOI21X1_1808 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_21_), .B(_12711_), .C(_12773_), .Y(_12721_) );
NOR2X1 NOR2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf0), .B(nonce_iniciales[85]), .Y(_12722_) );
AOI21X1 AOI21X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_12721_), .B(_12720_), .C(_12722_), .Y(_12592__21_) );
NOR2X1 NOR2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_12716_), .B(_12712_), .Y(_12723_) );
INVX1 INVX1_1785 ( .gnd(gnd), .vdd(vdd), .A(_12723_), .Y(_12724_) );
OAI21X1 OAI21X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_12718_), .B(_12724_), .C(module_2_W_22_), .Y(_12725_) );
INVX1 INVX1_1786 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_22_), .Y(_12726_) );
NAND3X1 NAND3X1_2922 ( .gnd(gnd), .vdd(vdd), .A(_12726_), .B(_12723_), .C(_12710_), .Y(_12727_) );
AND2X2 AND2X2_284 ( .gnd(gnd), .vdd(vdd), .A(_12725_), .B(_12727_), .Y(_12728_) );
NOR2X1 NOR2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf0), .B(nonce_iniciales[86]), .Y(_12729_) );
AOI21X1 AOI21X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_12628__bF_buf3), .B(_12728_), .C(_12729_), .Y(_12592__22_) );
NOR2X1 NOR2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf1), .B(nonce_iniciales[87]), .Y(_12730_) );
INVX1 INVX1_1787 ( .gnd(gnd), .vdd(vdd), .A(_12616_), .Y(_12731_) );
NAND3X1 NAND3X1_2923 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_20_), .B(_12731_), .C(_12710_), .Y(_12732_) );
OR2X2 OR2X2_302 ( .gnd(gnd), .vdd(vdd), .A(_12732_), .B(module_2_W_23_), .Y(_12733_) );
AOI21X1 AOI21X1_1811 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_23_), .B(_12732_), .C(_12665_), .Y(_12734_) );
AOI21X1 AOI21X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_12733_), .B(_12734_), .C(_12730_), .Y(_12592__23_) );
NOR2X1 NOR2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_12619_), .B(_12696_), .Y(_12735_) );
XNOR2X1 XNOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_12735_), .B(module_2_W_24_), .Y(_12736_) );
NOR2X1 NOR2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf1), .B(nonce_iniciales[88]), .Y(_12737_) );
AOI21X1 AOI21X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_12628__bF_buf3), .B(_12736_), .C(_12737_), .Y(_12592__24_) );
INVX1 INVX1_1788 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_25_), .Y(_12738_) );
AND2X2 AND2X2_285 ( .gnd(gnd), .vdd(vdd), .A(_12735_), .B(module_2_W_24_), .Y(_12739_) );
AOI21X1 AOI21X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_12738_), .B(_12739_), .C(_12717_), .Y(_12740_) );
NAND2X1 NAND2X1_1710 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_24_), .B(_12735_), .Y(_12741_) );
AOI21X1 AOI21X1_1815 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_25_), .B(_12741_), .C(_12773_), .Y(_12742_) );
NOR2X1 NOR2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf1), .B(nonce_iniciales[89]), .Y(_12743_) );
AOI21X1 AOI21X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_12742_), .B(_12740_), .C(_12743_), .Y(_12592__25_) );
NOR3X1 NOR3X1_374 ( .gnd(gnd), .vdd(vdd), .A(_12599_), .B(_12619_), .C(_12696_), .Y(_12744_) );
XNOR2X1 XNOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_12744_), .B(module_2_W_26_), .Y(_12745_) );
NOR2X1 NOR2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf1), .B(nonce_iniciales[90]), .Y(_12746_) );
AOI21X1 AOI21X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_12628__bF_buf3), .B(_12745_), .C(_12746_), .Y(_12592__26_) );
NOR2X1 NOR2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf1), .B(nonce_iniciales[91]), .Y(_12747_) );
AND2X2 AND2X2_286 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_26_), .B(module_2_W_25_), .Y(_12748_) );
NAND3X1 NAND3X1_2924 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_24_), .B(_12748_), .C(_12735_), .Y(_12749_) );
OR2X2 OR2X2_303 ( .gnd(gnd), .vdd(vdd), .A(_12749_), .B(module_2_W_27_), .Y(_12750_) );
AOI21X1 AOI21X1_1818 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_27_), .B(_12749_), .C(_12665_), .Y(_12751_) );
AOI21X1 AOI21X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_12750_), .B(_12751_), .C(_12747_), .Y(_12592__27_) );
INVX1 INVX1_1789 ( .gnd(gnd), .vdd(vdd), .A(_12601_), .Y(_12752_) );
NOR3X1 NOR3X1_375 ( .gnd(gnd), .vdd(vdd), .A(_12752_), .B(_12619_), .C(_12696_), .Y(_12753_) );
NAND2X1 NAND2X1_1711 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_28_), .B(_12753_), .Y(_12754_) );
INVX1 INVX1_1790 ( .gnd(gnd), .vdd(vdd), .A(_12619_), .Y(_12755_) );
NAND3X1 NAND3X1_2925 ( .gnd(gnd), .vdd(vdd), .A(_12601_), .B(_12755_), .C(_12690_), .Y(_12756_) );
NAND2X1 NAND2X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_12606_), .B(_12756_), .Y(_12757_) );
NAND2X1 NAND2X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_12754_), .B(_12757_), .Y(_12758_) );
NOR2X1 NOR2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf0), .B(nonce_iniciales[92]), .Y(_12759_) );
AOI21X1 AOI21X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_12628__bF_buf0), .B(_12758_), .C(_12759_), .Y(_12592__28_) );
NOR2X1 NOR2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf0), .B(nonce_iniciales[93]), .Y(_12760_) );
OR2X2 OR2X2_304 ( .gnd(gnd), .vdd(vdd), .A(_12754_), .B(module_2_W_29_), .Y(_12761_) );
AOI21X1 AOI21X1_1821 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_29_), .B(_12754_), .C(_12665_), .Y(_12762_) );
AOI21X1 AOI21X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_12761_), .B(_12762_), .C(_12760_), .Y(_12592__29_) );
NAND3X1 NAND3X1_2926 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_30_), .B(_12607_), .C(_12753_), .Y(_12763_) );
INVX1 INVX1_1791 ( .gnd(gnd), .vdd(vdd), .A(_12607_), .Y(_12764_) );
OAI21X1 OAI21X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_12756_), .B(_12764_), .C(_12609_), .Y(_12765_) );
NAND2X1 NAND2X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_12763_), .B(_12765_), .Y(_12766_) );
NOR2X1 NOR2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf8), .B(nonce_iniciales[94]), .Y(_12767_) );
AOI21X1 AOI21X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_12628__bF_buf0), .B(_12766_), .C(_12767_), .Y(_12592__30_) );
NOR2X1 NOR2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf0), .B(nonce_iniciales[95]), .Y(_12768_) );
NOR2X1 NOR2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_12764_), .B(_12756_), .Y(_12769_) );
NAND3X1 NAND3X1_2927 ( .gnd(gnd), .vdd(vdd), .A(_12608_), .B(module_2_W_30_), .C(_12769_), .Y(_12770_) );
AOI21X1 AOI21X1_1824 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_31_), .B(_12763_), .C(_12665_), .Y(_12771_) );
AOI21X1 AOI21X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_12770_), .B(_12771_), .C(_12768_), .Y(_12592__31_) );
DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__0_), .Q(module_2_W_0_) );
DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__1_), .Q(module_2_W_1_) );
DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__2_), .Q(module_2_W_2_) );
DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__3_), .Q(module_2_W_3_) );
DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__4_), .Q(module_2_W_4_) );
DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__5_), .Q(module_2_W_5_) );
DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__6_), .Q(module_2_W_6_) );
DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__7_), .Q(module_2_W_7_) );
DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__8_), .Q(module_2_W_8_) );
DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__9_), .Q(module_2_W_9_) );
DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__10_), .Q(module_2_W_10_) );
DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__11_), .Q(module_2_W_11_) );
DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__12_), .Q(module_2_W_12_) );
DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__13_), .Q(module_2_W_13_) );
DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__14_), .Q(module_2_W_14_) );
DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12592__15_), .Q(module_2_W_15_) );
DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__16_), .Q(module_2_W_16_) );
DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_12592__17_), .Q(module_2_W_17_) );
DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_12592__18_), .Q(module_2_W_18_) );
DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_12592__19_), .Q(module_2_W_19_) );
DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_12592__20_), .Q(module_2_W_20_) );
DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__21_), .Q(module_2_W_21_) );
DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__22_), .Q(module_2_W_22_) );
DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_12592__23_), .Q(module_2_W_23_) );
DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_12592__24_), .Q(module_2_W_24_) );
DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_12592__25_), .Q(module_2_W_25_) );
DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__26_), .Q(module_2_W_26_) );
DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_12592__27_), .Q(module_2_W_27_) );
DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__28_), .Q(module_2_W_28_) );
DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__29_), .Q(module_2_W_29_) );
DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__30_), .Q(module_2_W_30_) );
DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12592__31_), .Q(module_2_W_31_) );
INVX1 INVX1_1792 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_12811_) );
INVX1 INVX1_1793 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .Y(_12812_) );
INVX1 INVX1_1794 ( .gnd(gnd), .vdd(vdd), .A(target[0]), .Y(_12813_) );
OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_12812_), .B(gnd), .C(_12813_), .D(vdd), .Y(_12814_) );
OAI21X1 OAI21X1_2051 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .B(_12811_), .C(_12814_), .Y(_12815_) );
XOR2X1 XOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(vdd), .Y(_12816_) );
INVX2 INVX2_447 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .Y(_12817_) );
INVX1 INVX1_1795 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_12818_) );
NAND2X1 NAND2X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_12817_), .B(_12818_), .Y(_12819_) );
NAND2X1 NAND2X1_1716 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(gnd), .Y(_12820_) );
AOI21X1 AOI21X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_12819_), .B(_12820_), .C(_12816_), .Y(_12821_) );
INVX1 INVX1_1796 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .Y(_12822_) );
NAND2X1 NAND2X1_1717 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_12822_), .Y(_12823_) );
NAND2X1 NAND2X1_1718 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_12817_), .Y(_12824_) );
OAI21X1 OAI21X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_12816_), .B(_12824_), .C(_12823_), .Y(_12825_) );
AOI21X1 AOI21X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_12815_), .B(_12821_), .C(_12825_), .Y(_12826_) );
INVX1 INVX1_1797 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_15_), .Y(_12827_) );
INVX1 INVX1_1798 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_14_), .Y(_12828_) );
OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_12827_), .B(target[7]), .C(target[6]), .D(_12828_), .Y(_12829_) );
INVX4 INVX4_12 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .Y(_12830_) );
INVX2 INVX2_448 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .Y(_12831_) );
OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_12830_), .B(module_2_H_15_), .C(_12831_), .D(module_2_H_14_), .Y(_12832_) );
NOR2X1 NOR2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_12829_), .B(_12832_), .Y(_12833_) );
INVX2 INVX2_449 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_13_), .Y(_12834_) );
INVX1 INVX1_1799 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_12_), .Y(_12835_) );
OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_12834_), .B(target[5]), .C(target[4]), .D(_12835_), .Y(_12836_) );
INVX2 INVX2_450 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .Y(_12837_) );
INVX1 INVX1_1800 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .Y(_12838_) );
OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_12837_), .B(module_2_H_13_), .C(_12838_), .D(module_2_H_12_), .Y(_12839_) );
NOR2X1 NOR2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_12836_), .B(_12839_), .Y(_12840_) );
NAND2X1 NAND2X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_12833_), .B(_12840_), .Y(_12841_) );
NAND2X1 NAND2X1_1720 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .B(_12834_), .Y(_12842_) );
NAND3X1 NAND3X1_2928 ( .gnd(gnd), .vdd(vdd), .A(_12836_), .B(_12842_), .C(_12833_), .Y(_12843_) );
OAI21X1 OAI21X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_12826_), .B(_12841_), .C(_12843_), .Y(_12844_) );
INVX1 INVX1_1801 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_17_), .Y(_12845_) );
OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_12812_), .B(module_2_H_17_), .C(_12813_), .D(module_2_H_16_), .Y(_12846_) );
OAI21X1 OAI21X1_2054 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .B(_12845_), .C(_12846_), .Y(_12847_) );
XOR2X1 XOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(module_2_H_19_), .Y(_12848_) );
INVX1 INVX1_1802 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_18_), .Y(_12849_) );
NAND2X1 NAND2X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_12817_), .B(_12849_), .Y(_12850_) );
NAND2X1 NAND2X1_1722 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(module_2_H_18_), .Y(_12851_) );
AOI21X1 AOI21X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_12850_), .B(_12851_), .C(_12848_), .Y(_12852_) );
NAND2X1 NAND2X1_1723 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_19_), .B(_12822_), .Y(_12774_) );
NAND2X1 NAND2X1_1724 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_18_), .B(_12817_), .Y(_12775_) );
OAI21X1 OAI21X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_12848_), .B(_12775_), .C(_12774_), .Y(_12776_) );
AOI21X1 AOI21X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_12847_), .B(_12852_), .C(_12776_), .Y(_12777_) );
INVX1 INVX1_1803 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_23_), .Y(_12778_) );
INVX1 INVX1_1804 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_22_), .Y(_12779_) );
OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_12778_), .B(target[7]), .C(target[6]), .D(_12779_), .Y(_12780_) );
OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_12830_), .B(module_2_H_23_), .C(_12831_), .D(module_2_H_22_), .Y(_12781_) );
NOR2X1 NOR2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_12781_), .Y(_12782_) );
NAND2X1 NAND2X1_1725 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_21_), .B(_12837_), .Y(_12783_) );
NAND2X1 NAND2X1_1726 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_20_), .B(_12838_), .Y(_12784_) );
AND2X2 AND2X2_287 ( .gnd(gnd), .vdd(vdd), .A(_12783_), .B(_12784_), .Y(_12785_) );
INVX1 INVX1_1805 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_20_), .Y(_12786_) );
NOR2X1 NOR2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_21_), .B(_12837_), .Y(_12787_) );
AOI21X1 AOI21X1_1830 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_12786_), .C(_12787_), .Y(_12788_) );
NAND3X1 NAND3X1_2929 ( .gnd(gnd), .vdd(vdd), .A(_12785_), .B(_12788_), .C(_12782_), .Y(_12789_) );
AOI21X1 AOI21X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_12783_), .B(_12784_), .C(_12787_), .Y(_12790_) );
AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_12830_), .B(module_2_H_23_), .C(_12831_), .D(module_2_H_22_), .Y(_12791_) );
NOR2X1 NOR2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_23_), .B(_12830_), .Y(_12792_) );
AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_12830_), .B(module_2_H_15_), .C(_12831_), .D(module_2_H_14_), .Y(_12793_) );
NOR2X1 NOR2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_15_), .B(_12830_), .Y(_12794_) );
OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_12791_), .B(_12792_), .C(_12793_), .D(_12794_), .Y(_12795_) );
AOI21X1 AOI21X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_12782_), .B(_12790_), .C(_12795_), .Y(_12796_) );
OAI21X1 OAI21X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_12777_), .B(_12789_), .C(_12796_), .Y(_12797_) );
NOR2X1 NOR2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf3), .B(_12797__bF_buf3), .Y(module_2_comparador_target_hash_0_terminado) );
INVX1 INVX1_1806 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_0_), .Y(_12798_) );
NOR3X1 NOR3X1_376 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf0), .B(_12798_), .C(_12797__bF_buf0), .Y(bounty_48_) );
INVX1 INVX1_1807 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_1_), .Y(_12799_) );
NOR3X1 NOR3X1_377 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf4), .B(_12799_), .C(_12797__bF_buf2), .Y(bounty_49_) );
INVX1 INVX1_1808 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_2_), .Y(_12800_) );
NOR3X1 NOR3X1_378 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf4), .B(_12800_), .C(_12797__bF_buf2), .Y(bounty_50_) );
INVX1 INVX1_1809 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_3_), .Y(_12801_) );
NOR3X1 NOR3X1_379 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf2), .B(_12801_), .C(_12797__bF_buf4), .Y(bounty_51_) );
INVX1 INVX1_1810 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_4_), .Y(_12802_) );
NOR3X1 NOR3X1_380 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf4), .B(_12802_), .C(_12797__bF_buf2), .Y(bounty_52_) );
INVX1 INVX1_1811 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_5_), .Y(_12803_) );
NOR3X1 NOR3X1_381 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf2), .B(_12803_), .C(_12797__bF_buf4), .Y(bounty_53_) );
INVX1 INVX1_1812 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_6_), .Y(_12804_) );
NOR3X1 NOR3X1_382 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf2), .B(_12804_), .C(_12797__bF_buf4), .Y(bounty_54_) );
INVX1 INVX1_1813 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_7_), .Y(_12805_) );
NOR3X1 NOR3X1_383 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf2), .B(_12805_), .C(_12797__bF_buf4), .Y(bounty_55_) );
INVX1 INVX1_1814 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_12806_) );
NOR3X1 NOR3X1_384 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf3), .B(_12806_), .C(_12797__bF_buf3), .Y(bounty_56_) );
NOR3X1 NOR3X1_385 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf3), .B(_12811_), .C(_12797__bF_buf3), .Y(bounty_57_) );
NOR3X1 NOR3X1_386 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf1), .B(_12818_), .C(_12797__bF_buf1), .Y(bounty_58_) );
INVX1 INVX1_1815 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_12807_) );
NOR3X1 NOR3X1_387 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf3), .B(_12807_), .C(_12797__bF_buf3), .Y(bounty_59_) );
NOR3X1 NOR3X1_388 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf0), .B(_12835_), .C(_12797__bF_buf0), .Y(bounty_60_) );
NOR3X1 NOR3X1_389 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf2), .B(_12834_), .C(_12797__bF_buf4), .Y(bounty_61_) );
NOR3X1 NOR3X1_390 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf4), .B(_12828_), .C(_12797__bF_buf2), .Y(bounty_62_) );
NOR3X1 NOR3X1_391 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf4), .B(_12827_), .C(_12797__bF_buf2), .Y(bounty_63_) );
INVX1 INVX1_1816 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_16_), .Y(_12808_) );
NOR3X1 NOR3X1_392 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf3), .B(_12808_), .C(_12797__bF_buf3), .Y(bounty_64_) );
NOR3X1 NOR3X1_393 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf1), .B(_12845_), .C(_12797__bF_buf1), .Y(bounty_65_) );
NOR3X1 NOR3X1_394 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf1), .B(_12849_), .C(_12797__bF_buf1), .Y(bounty_66_) );
INVX1 INVX1_1817 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_19_), .Y(_12809_) );
NOR3X1 NOR3X1_395 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf1), .B(_12809_), .C(_12797__bF_buf1), .Y(bounty_67_) );
NOR3X1 NOR3X1_396 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf0), .B(_12786_), .C(_12797__bF_buf0), .Y(bounty_68_) );
INVX1 INVX1_1818 ( .gnd(gnd), .vdd(vdd), .A(module_2_H_21_), .Y(_12810_) );
NOR3X1 NOR3X1_397 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf1), .B(_12810_), .C(_12797__bF_buf1), .Y(bounty_69_) );
NOR3X1 NOR3X1_398 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf0), .B(_12779_), .C(_12797__bF_buf0), .Y(bounty_70_) );
NOR3X1 NOR3X1_399 ( .gnd(gnd), .vdd(vdd), .A(_12844__bF_buf0), .B(_12778_), .C(_12797__bF_buf0), .Y(bounty_71_) );
INVX1 INVX1_1819 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf4_), .Y(_12853_) );
AOI21X1 AOI21X1_1833 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_24_), .B(_12853_), .C(bloque_datos_80_bF_buf4_), .Y(_12854_) );
OAI21X1 OAI21X1_2057 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_24_), .B(_12853_), .C(_12854_), .Y(module_2_W_136_) );
INVX1 INVX1_1820 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf0_), .Y(_12855_) );
AOI21X1 AOI21X1_1834 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_25_), .B(_12855_), .C(bloque_datos_81_bF_buf0_), .Y(_12856_) );
OAI21X1 OAI21X1_2058 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_25_), .B(_12855_), .C(_12856_), .Y(module_2_W_137_) );
INVX1 INVX1_1821 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf4_), .Y(_12857_) );
AOI21X1 AOI21X1_1835 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_26_), .B(_12857_), .C(bloque_datos_82_bF_buf3_), .Y(_12858_) );
OAI21X1 OAI21X1_2059 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_26_), .B(_12857_), .C(_12858_), .Y(module_2_W_138_) );
INVX1 INVX1_1822 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf4_), .Y(_12859_) );
AOI21X1 AOI21X1_1836 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_27_), .B(_12859_), .C(bloque_datos_83_bF_buf4_), .Y(_12860_) );
OAI21X1 OAI21X1_2060 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_27_), .B(_12859_), .C(_12860_), .Y(module_2_W_139_) );
INVX1 INVX1_1823 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf2_), .Y(_12861_) );
AOI21X1 AOI21X1_1837 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_28_), .B(_12861_), .C(bloque_datos_84_bF_buf4_), .Y(_12862_) );
OAI21X1 OAI21X1_2061 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_28_), .B(_12861_), .C(_12862_), .Y(module_2_W_140_) );
INVX1 INVX1_1824 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf2_), .Y(_12863_) );
AOI21X1 AOI21X1_1838 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_29_), .B(_12863_), .C(bloque_datos_85_bF_buf2_), .Y(_12864_) );
OAI21X1 OAI21X1_2062 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_29_), .B(_12863_), .C(_12864_), .Y(module_2_W_141_) );
INVX1 INVX1_1825 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf2_), .Y(_12865_) );
AOI21X1 AOI21X1_1839 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_30_), .B(_12865_), .C(bloque_datos_86_bF_buf4_), .Y(_12866_) );
OAI21X1 OAI21X1_2063 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_30_), .B(_12865_), .C(_12866_), .Y(module_2_W_142_) );
INVX1 INVX1_1826 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .Y(_12867_) );
AOI21X1 AOI21X1_1840 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_31_), .B(_12867_), .C(bloque_datos_87_bF_buf3_), .Y(_12868_) );
OAI21X1 OAI21X1_2064 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_31_), .B(_12867_), .C(_12868_), .Y(module_2_W_143_) );
INVX1 INVX1_1827 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf0_), .Y(_12869_) );
OR2X2 OR2X2_305 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_16_), .B(bloque_datos_24_bF_buf4_), .Y(_12870_) );
NAND2X1 NAND2X1_1727 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_16_), .B(bloque_datos_24_bF_buf3_), .Y(_12871_) );
NAND2X1 NAND2X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_12871_), .B(_12870_), .Y(_12872_) );
NAND2X1 NAND2X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_12869_), .B(_12872_), .Y(module_2_W_128_) );
INVX1 INVX1_1828 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf3_), .Y(_12873_) );
AOI21X1 AOI21X1_1841 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_17_), .B(_12873_), .C(bloque_datos_73_bF_buf2_), .Y(_12874_) );
OAI21X1 OAI21X1_2065 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_17_), .B(_12873_), .C(_12874_), .Y(module_2_W_129_) );
INVX1 INVX1_1829 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf0_), .Y(_12875_) );
OR2X2 OR2X2_306 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_18_), .B(bloque_datos_26_bF_buf2_), .Y(_12876_) );
NAND2X1 NAND2X1_1730 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_18_), .B(bloque_datos_26_bF_buf1_), .Y(_12877_) );
NAND2X1 NAND2X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_12877_), .B(_12876_), .Y(_12878_) );
NAND2X1 NAND2X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_12875_), .B(_12878_), .Y(module_2_W_130_) );
INVX1 INVX1_1830 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf2_), .Y(_12879_) );
OR2X2 OR2X2_307 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_19_), .B(bloque_datos_27_bF_buf2_), .Y(_12880_) );
NAND2X1 NAND2X1_1733 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_19_), .B(bloque_datos_27_bF_buf1_), .Y(_12881_) );
NAND2X1 NAND2X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_12881_), .B(_12880_), .Y(_12882_) );
NAND2X1 NAND2X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_12879_), .B(_12882_), .Y(module_2_W_131_) );
INVX2 INVX2_451 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf2_), .Y(_12883_) );
AOI21X1 AOI21X1_1842 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_20_), .B(_12883_), .C(bloque_datos_76_bF_buf4_), .Y(_12884_) );
OAI21X1 OAI21X1_2066 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_20_), .B(_12883_), .C(_12884_), .Y(module_2_W_132_) );
INVX2 INVX2_452 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf2_), .Y(_12885_) );
AOI21X1 AOI21X1_1843 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_21_), .B(_12885_), .C(bloque_datos_77_bF_buf4_), .Y(_12886_) );
OAI21X1 OAI21X1_2067 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_21_), .B(_12885_), .C(_12886_), .Y(module_2_W_133_) );
INVX2 INVX2_453 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf2_), .Y(_12887_) );
AOI21X1 AOI21X1_1844 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_22_), .B(_12887_), .C(bloque_datos_78_bF_buf4_), .Y(_12888_) );
OAI21X1 OAI21X1_2068 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_22_), .B(_12887_), .C(_12888_), .Y(module_2_W_134_) );
INVX1 INVX1_1831 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf1_), .Y(_12889_) );
AOI21X1 AOI21X1_1845 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_23_), .B(_12889_), .C(bloque_datos_79_bF_buf2_), .Y(_12890_) );
OAI21X1 OAI21X1_2069 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_23_), .B(_12889_), .C(_12890_), .Y(module_2_W_135_) );
INVX1 INVX1_1832 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(_12891_) );
INVX1 INVX1_1833 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf2_), .Y(_12892_) );
OAI21X1 OAI21X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_12891_), .B(bloque_datos_40_bF_buf4_), .C(_12892_), .Y(_12893_) );
AOI21X1 AOI21X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_12891_), .B(bloque_datos_40_bF_buf3_), .C(_12893_), .Y(_12894_) );
INVX1 INVX1_1834 ( .gnd(gnd), .vdd(vdd), .A(_12894_), .Y(module_2_W_144_) );
INVX1 INVX1_1835 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(_12895_) );
INVX1 INVX1_1836 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf0_), .Y(_12896_) );
OAI21X1 OAI21X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_12895_), .B(bloque_datos_41_bF_buf3_), .C(_12896_), .Y(_12897_) );
AOI21X1 AOI21X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_12895_), .B(bloque_datos_41_bF_buf2_), .C(_12897_), .Y(_12898_) );
INVX1 INVX1_1837 ( .gnd(gnd), .vdd(vdd), .A(_12898_), .Y(module_2_W_145_) );
INVX1 INVX1_1838 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf0_), .Y(_12899_) );
INVX1 INVX1_1839 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf2_), .Y(_12900_) );
OAI21X1 OAI21X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_12899_), .B(bloque_datos_42_bF_buf3_), .C(_12900_), .Y(_12901_) );
AOI21X1 AOI21X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_12899_), .B(bloque_datos_42_bF_buf2_), .C(_12901_), .Y(_12902_) );
INVX1 INVX1_1840 ( .gnd(gnd), .vdd(vdd), .A(_12902_), .Y(module_2_W_146_) );
INVX1 INVX1_1841 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf0_), .Y(_12903_) );
INVX1 INVX1_1842 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf2_), .Y(_12904_) );
OAI21X1 OAI21X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_12903_), .B(bloque_datos_43_bF_buf3_), .C(_12904_), .Y(_12905_) );
AOI21X1 AOI21X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_12903_), .B(bloque_datos_43_bF_buf2_), .C(_12905_), .Y(_12906_) );
INVX1 INVX1_1843 ( .gnd(gnd), .vdd(vdd), .A(_12906_), .Y(module_2_W_147_) );
INVX1 INVX1_1844 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf0_), .Y(_12907_) );
INVX1 INVX1_1845 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf0_), .Y(_12908_) );
OAI21X1 OAI21X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_12907_), .B(bloque_datos_44_bF_buf4_), .C(_12908_), .Y(_12909_) );
AOI21X1 AOI21X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_12907_), .B(bloque_datos_44_bF_buf3_), .C(_12909_), .Y(_12910_) );
INVX1 INVX1_1846 ( .gnd(gnd), .vdd(vdd), .A(_12910_), .Y(module_2_W_148_) );
INVX1 INVX1_1847 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf0_), .Y(_12911_) );
INVX1 INVX1_1848 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf0_), .Y(_12912_) );
OAI21X1 OAI21X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_12911_), .B(bloque_datos_45_bF_buf4_), .C(_12912_), .Y(_12913_) );
AOI21X1 AOI21X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_12911_), .B(bloque_datos_45_bF_buf3_), .C(_12913_), .Y(_12914_) );
INVX1 INVX1_1849 ( .gnd(gnd), .vdd(vdd), .A(_12914_), .Y(module_2_W_149_) );
INVX1 INVX1_1850 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf0_), .Y(_12915_) );
INVX1 INVX1_1851 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf0_), .Y(_12916_) );
OAI21X1 OAI21X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_12915_), .B(bloque_datos_46_bF_buf4_), .C(_12916_), .Y(_12917_) );
AOI21X1 AOI21X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_12915_), .B(bloque_datos_46_bF_buf3_), .C(_12917_), .Y(_12918_) );
INVX2 INVX2_454 ( .gnd(gnd), .vdd(vdd), .A(_12918_), .Y(module_2_W_150_) );
INVX1 INVX1_1852 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[7]), .Y(_12919_) );
INVX1 INVX1_1853 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf1_), .Y(_12920_) );
OAI21X1 OAI21X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_12919_), .B(bloque_datos_47_bF_buf2_), .C(_12920_), .Y(_12921_) );
AOI21X1 AOI21X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_12919_), .B(bloque_datos_47_bF_buf1_), .C(_12921_), .Y(_12922_) );
INVX2 INVX2_455 ( .gnd(gnd), .vdd(vdd), .A(_12922_), .Y(module_2_W_151_) );
AOI21X1 AOI21X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_12871_), .B(_12870_), .C(bloque_datos_72_bF_buf4_), .Y(_12923_) );
XNOR2X1 XNOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .B(bloque_datos_48_bF_buf4_), .Y(_12924_) );
NAND2X1 NAND2X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_12924_), .B(_12923_), .Y(module_2_W_152_) );
XOR2X1 XOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .B(bloque_datos_49_bF_buf2_), .Y(_12925_) );
NOR2X1 NOR2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_12925_), .B(module_2_W_129_), .Y(_12926_) );
INVX1 INVX1_1854 ( .gnd(gnd), .vdd(vdd), .A(_12926_), .Y(module_2_W_153_) );
AOI21X1 AOI21X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_12877_), .B(_12876_), .C(bloque_datos_74_bF_buf4_), .Y(_12927_) );
XNOR2X1 XNOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .B(bloque_datos_50_bF_buf3_), .Y(_12928_) );
NAND2X1 NAND2X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_12928_), .B(_12927_), .Y(module_2_W_154_) );
AOI21X1 AOI21X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_12881_), .B(_12880_), .C(bloque_datos_75_bF_buf1_), .Y(_12929_) );
XNOR2X1 XNOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .B(bloque_datos_51_bF_buf3_), .Y(_12930_) );
NAND2X1 NAND2X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_12930_), .B(_12929_), .Y(module_2_W_155_) );
INVX1 INVX1_1855 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_20_), .Y(_12931_) );
INVX1 INVX1_1856 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf3_), .Y(_12932_) );
OAI21X1 OAI21X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_12931_), .B(bloque_datos_28_bF_buf1_), .C(_12932_), .Y(_12933_) );
AOI21X1 AOI21X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_12931_), .B(bloque_datos_28_bF_buf0_), .C(_12933_), .Y(_12934_) );
AND2X2 AND2X2_288 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf2_), .B(bloque_datos_52_bF_buf4_), .Y(_12935_) );
NOR2X1 NOR2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf1_), .B(bloque_datos_52_bF_buf3_), .Y(_12936_) );
OAI21X1 OAI21X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_12935_), .B(_12936_), .C(_12934_), .Y(module_2_W_156_) );
XOR2X1 XOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf0_), .B(bloque_datos_53_bF_buf2_), .Y(_12937_) );
NOR2X1 NOR2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_12937_), .B(module_2_W_133_), .Y(_12938_) );
INVX1 INVX1_1857 ( .gnd(gnd), .vdd(vdd), .A(_12938_), .Y(module_2_W_157_) );
XOR2X1 XOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf0_), .B(bloque_datos_54_bF_buf2_), .Y(_12939_) );
NOR2X1 NOR2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_12939_), .B(module_2_W_134_), .Y(_12940_) );
INVX1 INVX1_1858 ( .gnd(gnd), .vdd(vdd), .A(_12940_), .Y(module_2_W_158_) );
XOR2X1 XOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[15]), .B(bloque_datos[55]), .Y(_12941_) );
NOR2X1 NOR2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_12941_), .B(module_2_W_135_), .Y(_12942_) );
INVX1 INVX1_1859 ( .gnd(gnd), .vdd(vdd), .A(_12942_), .Y(module_2_W_159_) );
XOR2X1 XOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_24_), .B(bloque_datos_32_bF_buf3_), .Y(_12943_) );
NOR2X1 NOR2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf3_), .B(_12943_), .Y(_12944_) );
XNOR2X1 XNOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf0_), .B(bloque_datos_56_bF_buf4_), .Y(_12945_) );
NAND2X1 NAND2X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_12945_), .B(_12944_), .Y(module_2_W_160_) );
INVX1 INVX1_1860 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_25_), .Y(_12946_) );
INVX1 INVX1_1861 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf4_), .Y(_12947_) );
OAI21X1 OAI21X1_2080 ( .gnd(gnd), .vdd(vdd), .A(_12946_), .B(bloque_datos_33_bF_buf3_), .C(_12947_), .Y(_12948_) );
AOI21X1 AOI21X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_12946_), .B(bloque_datos_33_bF_buf2_), .C(_12948_), .Y(_12949_) );
XNOR2X1 XNOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .B(bloque_datos_57_bF_buf3_), .Y(_12950_) );
NAND2X1 NAND2X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_12950_), .B(_12949_), .Y(module_2_W_161_) );
XOR2X1 XOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_26_), .B(bloque_datos_34_bF_buf3_), .Y(_12951_) );
NOR2X1 NOR2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf2_), .B(_12951_), .Y(_12952_) );
XNOR2X1 XNOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .B(bloque_datos_58_bF_buf4_), .Y(_12953_) );
NAND2X1 NAND2X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_12953_), .B(_12952_), .Y(module_2_W_162_) );
XOR2X1 XOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_27_), .B(bloque_datos_35_bF_buf3_), .Y(_12954_) );
NOR2X1 NOR2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf3_), .B(_12954_), .Y(_12955_) );
XNOR2X1 XNOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf0_), .B(bloque_datos_59_bF_buf4_), .Y(_12956_) );
NAND2X1 NAND2X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_12956_), .B(_12955_), .Y(module_2_W_163_) );
XOR2X1 XOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf0_), .B(bloque_datos_60_bF_buf2_), .Y(_12957_) );
NOR2X1 NOR2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_12957_), .B(module_2_W_140_), .Y(_12958_) );
INVX1 INVX1_1862 ( .gnd(gnd), .vdd(vdd), .A(_12958_), .Y(module_2_W_164_) );
XOR2X1 XOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf0_), .B(bloque_datos_61_bF_buf4_), .Y(_12959_) );
NOR2X1 NOR2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_12959_), .B(module_2_W_141_), .Y(_12960_) );
INVX1 INVX1_1863 ( .gnd(gnd), .vdd(vdd), .A(_12960_), .Y(module_2_W_165_) );
XOR2X1 XOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf0_), .B(bloque_datos_62_bF_buf2_), .Y(_12961_) );
NOR2X1 NOR2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_12961_), .B(module_2_W_142_), .Y(_12962_) );
INVX2 INVX2_456 ( .gnd(gnd), .vdd(vdd), .A(_12962_), .Y(module_2_W_166_) );
XOR2X1 XOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf0_), .B(bloque_datos[63]), .Y(_12963_) );
NOR2X1 NOR2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_12963_), .B(module_2_W_143_), .Y(_12964_) );
INVX1 INVX1_1864 ( .gnd(gnd), .vdd(vdd), .A(_12964_), .Y(module_2_W_167_) );
XNOR2X1 XNOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf2_), .B(bloque_datos_64_bF_buf4_), .Y(_12965_) );
AND2X2 AND2X2_289 ( .gnd(gnd), .vdd(vdd), .A(_12894_), .B(_12965_), .Y(_12966_) );
INVX2 INVX2_457 ( .gnd(gnd), .vdd(vdd), .A(_12966_), .Y(module_2_W_168_) );
XNOR2X1 XNOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf2_), .B(bloque_datos_65_bF_buf3_), .Y(_12967_) );
AND2X2 AND2X2_290 ( .gnd(gnd), .vdd(vdd), .A(_12898_), .B(_12967_), .Y(_12968_) );
INVX1 INVX1_1865 ( .gnd(gnd), .vdd(vdd), .A(_12968_), .Y(module_2_W_169_) );
XNOR2X1 XNOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf0_), .B(bloque_datos_66_bF_buf4_), .Y(_12969_) );
AND2X2 AND2X2_291 ( .gnd(gnd), .vdd(vdd), .A(_12902_), .B(_12969_), .Y(_12970_) );
INVX1 INVX1_1866 ( .gnd(gnd), .vdd(vdd), .A(_12970_), .Y(module_2_W_170_) );
AND2X2 AND2X2_292 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf0_), .B(bloque_datos_67_bF_buf2_), .Y(_12971_) );
NOR2X1 NOR2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf4_), .B(bloque_datos_67_bF_buf1_), .Y(_12972_) );
OAI21X1 OAI21X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_12971_), .B(_12972_), .C(_12906_), .Y(module_2_W_171_) );
INVX2 INVX2_458 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf2_), .Y(_12973_) );
NOR2X1 NOR2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_12883_), .B(_12973_), .Y(_12974_) );
NOR2X1 NOR2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf4_), .B(bloque_datos_68_bF_buf1_), .Y(_12975_) );
OAI21X1 OAI21X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_12974_), .B(_12975_), .C(_12910_), .Y(module_2_W_172_) );
INVX2 INVX2_459 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf2_), .Y(_12976_) );
NOR2X1 NOR2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_12885_), .B(_12976_), .Y(_12977_) );
NOR2X1 NOR2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf1_), .B(bloque_datos_69_bF_buf1_), .Y(_12978_) );
OAI21X1 OAI21X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_12977_), .B(_12978_), .C(_12914_), .Y(module_2_W_173_) );
INVX2 INVX2_460 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf2_), .Y(_12979_) );
NOR2X1 NOR2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_12887_), .B(_12979_), .Y(_12980_) );
NOR2X1 NOR2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf1_), .B(bloque_datos_70_bF_buf1_), .Y(_12981_) );
OAI21X1 OAI21X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_12980_), .B(_12981_), .C(_12918_), .Y(module_2_W_174_) );
XNOR2X1 XNOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf0_), .B(bloque_datos_71_bF_buf1_), .Y(_12982_) );
AND2X2 AND2X2_293 ( .gnd(gnd), .vdd(vdd), .A(_12922_), .B(_12982_), .Y(_12983_) );
INVX1 INVX1_1867 ( .gnd(gnd), .vdd(vdd), .A(_12983_), .Y(module_2_W_175_) );
XNOR2X1 XNOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf2_), .B(bloque_datos_72_bF_buf3_), .Y(_12984_) );
NAND3X1 NAND3X1_2930 ( .gnd(gnd), .vdd(vdd), .A(_12924_), .B(_12984_), .C(_12923_), .Y(module_2_W_176_) );
INVX1 INVX1_1868 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_17_), .Y(_12985_) );
NAND2X1 NAND2X1_1743 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf1_), .B(_12985_), .Y(_12986_) );
AND2X2 AND2X2_294 ( .gnd(gnd), .vdd(vdd), .A(_12874_), .B(_12986_), .Y(_12987_) );
INVX1 INVX1_1869 ( .gnd(gnd), .vdd(vdd), .A(_12925_), .Y(_12988_) );
XNOR2X1 XNOR2X1_339 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf1_), .B(bloque_datos_73_bF_buf1_), .Y(_12989_) );
NAND3X1 NAND3X1_2931 ( .gnd(gnd), .vdd(vdd), .A(_12988_), .B(_12989_), .C(_12987_), .Y(module_2_W_177_) );
XNOR2X1 XNOR2X1_340 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf2_), .B(bloque_datos_74_bF_buf3_), .Y(_12990_) );
NAND3X1 NAND3X1_2932 ( .gnd(gnd), .vdd(vdd), .A(_12928_), .B(_12990_), .C(_12927_), .Y(module_2_W_178_) );
XNOR2X1 XNOR2X1_341 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf2_), .B(bloque_datos_75_bF_buf0_), .Y(_12991_) );
NAND3X1 NAND3X1_2933 ( .gnd(gnd), .vdd(vdd), .A(_12930_), .B(_12991_), .C(_12929_), .Y(module_2_W_179_) );
XOR2X1 XOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf1_), .B(bloque_datos_76_bF_buf2_), .Y(_12992_) );
NOR2X1 NOR2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_12992_), .B(module_2_W_156_), .Y(_12993_) );
INVX1 INVX1_1870 ( .gnd(gnd), .vdd(vdd), .A(_12993_), .Y(module_2_W_180_) );
INVX1 INVX1_1871 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_21_), .Y(_12994_) );
INVX1 INVX1_1872 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf3_), .Y(_12995_) );
OAI21X1 OAI21X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_12994_), .B(bloque_datos_29_bF_buf0_), .C(_12995_), .Y(_12996_) );
AOI21X1 AOI21X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_12994_), .B(bloque_datos_29_bF_buf4_), .C(_12996_), .Y(_12997_) );
INVX1 INVX1_1873 ( .gnd(gnd), .vdd(vdd), .A(_12937_), .Y(_12998_) );
XNOR2X1 XNOR2X1_342 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf1_), .B(bloque_datos_77_bF_buf2_), .Y(_12999_) );
NAND3X1 NAND3X1_2934 ( .gnd(gnd), .vdd(vdd), .A(_12998_), .B(_12999_), .C(_12997_), .Y(module_2_W_181_) );
XNOR2X1 XNOR2X1_343 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf1_), .B(bloque_datos_78_bF_buf3_), .Y(_13000_) );
AND2X2 AND2X2_295 ( .gnd(gnd), .vdd(vdd), .A(_12940_), .B(_13000_), .Y(_13001_) );
INVX2 INVX2_461 ( .gnd(gnd), .vdd(vdd), .A(_13001_), .Y(module_2_W_182_) );
XNOR2X1 XNOR2X1_344 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .B(bloque_datos_79_bF_buf1_), .Y(_13002_) );
AND2X2 AND2X2_296 ( .gnd(gnd), .vdd(vdd), .A(_12942_), .B(_13002_), .Y(_13003_) );
INVX2 INVX2_462 ( .gnd(gnd), .vdd(vdd), .A(_13003_), .Y(module_2_W_183_) );
XNOR2X1 XNOR2X1_345 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf2_), .B(bloque_datos_40_bF_buf2_), .Y(_13004_) );
NAND3X1 NAND3X1_2935 ( .gnd(gnd), .vdd(vdd), .A(_12945_), .B(_13004_), .C(_12944_), .Y(module_2_W_184_) );
XNOR2X1 XNOR2X1_346 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf3_), .B(bloque_datos_41_bF_buf1_), .Y(_13005_) );
NAND3X1 NAND3X1_2936 ( .gnd(gnd), .vdd(vdd), .A(_12950_), .B(_13005_), .C(_12949_), .Y(module_2_W_185_) );
XNOR2X1 XNOR2X1_347 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf1_), .B(bloque_datos_42_bF_buf1_), .Y(_13006_) );
NAND3X1 NAND3X1_2937 ( .gnd(gnd), .vdd(vdd), .A(_12953_), .B(_13006_), .C(_12952_), .Y(module_2_W_186_) );
XNOR2X1 XNOR2X1_348 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf2_), .B(bloque_datos_43_bF_buf1_), .Y(_13007_) );
NAND3X1 NAND3X1_2938 ( .gnd(gnd), .vdd(vdd), .A(_12956_), .B(_13007_), .C(_12955_), .Y(module_2_W_187_) );
XNOR2X1 XNOR2X1_349 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf3_), .B(bloque_datos_44_bF_buf2_), .Y(_13008_) );
AND2X2 AND2X2_297 ( .gnd(gnd), .vdd(vdd), .A(_12958_), .B(_13008_), .Y(_13009_) );
INVX1 INVX1_1874 ( .gnd(gnd), .vdd(vdd), .A(_13009_), .Y(module_2_W_188_) );
XNOR2X1 XNOR2X1_350 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf1_), .B(bloque_datos_45_bF_buf2_), .Y(_13010_) );
AND2X2 AND2X2_298 ( .gnd(gnd), .vdd(vdd), .A(_12960_), .B(_13010_), .Y(_13011_) );
INVX1 INVX1_1875 ( .gnd(gnd), .vdd(vdd), .A(_13011_), .Y(module_2_W_189_) );
XNOR2X1 XNOR2X1_351 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf3_), .B(bloque_datos_46_bF_buf2_), .Y(_13012_) );
AND2X2 AND2X2_299 ( .gnd(gnd), .vdd(vdd), .A(_12962_), .B(_13012_), .Y(_13013_) );
INVX1 INVX1_1876 ( .gnd(gnd), .vdd(vdd), .A(_13013_), .Y(module_2_W_190_) );
XNOR2X1 XNOR2X1_352 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf2_), .B(bloque_datos_47_bF_buf0_), .Y(_13014_) );
AND2X2 AND2X2_300 ( .gnd(gnd), .vdd(vdd), .A(_12964_), .B(_13014_), .Y(_13015_) );
INVX1 INVX1_1877 ( .gnd(gnd), .vdd(vdd), .A(_13015_), .Y(module_2_W_191_) );
AND2X2 AND2X2_301 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf1_), .B(bloque_datos_48_bF_buf3_), .Y(_13016_) );
NOR2X1 NOR2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf0_), .B(bloque_datos_48_bF_buf2_), .Y(_13017_) );
OAI21X1 OAI21X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_13016_), .B(_13017_), .C(_12966_), .Y(module_2_W_192_) );
AND2X2 AND2X2_302 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf3_), .B(bloque_datos_49_bF_buf1_), .Y(_13018_) );
NOR2X1 NOR2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf2_), .B(bloque_datos_49_bF_buf0_), .Y(_13019_) );
OAI21X1 OAI21X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_13018_), .B(_13019_), .C(_12968_), .Y(module_2_W_193_) );
AND2X2 AND2X2_303 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf1_), .B(bloque_datos_50_bF_buf2_), .Y(_13020_) );
NOR2X1 NOR2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf0_), .B(bloque_datos_50_bF_buf1_), .Y(_13021_) );
OAI21X1 OAI21X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_13020_), .B(_13021_), .C(_12970_), .Y(module_2_W_194_) );
OR2X2 OR2X2_308 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_171_), .B(bloque_datos_51_bF_buf2_), .Y(module_2_W_195_) );
NOR2X1 NOR2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf2_), .B(module_2_W_172_), .Y(_13022_) );
INVX1 INVX1_1878 ( .gnd(gnd), .vdd(vdd), .A(_13022_), .Y(module_2_W_196_) );
NOR2X1 NOR2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf1_), .B(module_2_W_173_), .Y(_13023_) );
INVX1 INVX1_1879 ( .gnd(gnd), .vdd(vdd), .A(_13023_), .Y(module_2_W_197_) );
OR2X2 OR2X2_309 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_174_), .B(bloque_datos_54_bF_buf1_), .Y(module_2_W_198_) );
XNOR2X1 XNOR2X1_353 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf0_), .B(bloque_datos[55]), .Y(_13024_) );
NAND2X1 NAND2X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_13024_), .B(_12983_), .Y(module_2_W_199_) );
NAND2X1 NAND2X1_1745 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf3_), .B(module_2_W_128_), .Y(_13025_) );
INVX1 INVX1_1880 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf2_), .Y(_13026_) );
NAND2X1 NAND2X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_13026_), .B(_12923_), .Y(_13027_) );
AOI21X1 AOI21X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_13027_), .B(_13025_), .C(module_2_W_176_), .Y(_13028_) );
INVX2 INVX2_463 ( .gnd(gnd), .vdd(vdd), .A(_13028_), .Y(module_2_W_200_) );
NAND2X1 NAND2X1_1747 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf2_), .B(module_2_W_129_), .Y(_13029_) );
OR2X2 OR2X2_310 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_129_), .B(bloque_datos_57_bF_buf1_), .Y(_13030_) );
AOI21X1 AOI21X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_13029_), .B(_13030_), .C(module_2_W_177_), .Y(_13031_) );
INVX1 INVX1_1881 ( .gnd(gnd), .vdd(vdd), .A(_13031_), .Y(module_2_W_201_) );
NAND2X1 NAND2X1_1748 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf3_), .B(module_2_W_130_), .Y(_13032_) );
INVX1 INVX1_1882 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf2_), .Y(_13033_) );
NAND2X1 NAND2X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_13033_), .B(_12927_), .Y(_13034_) );
AOI21X1 AOI21X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_13034_), .B(_13032_), .C(module_2_W_178_), .Y(_13035_) );
INVX1 INVX1_1883 ( .gnd(gnd), .vdd(vdd), .A(_13035_), .Y(module_2_W_202_) );
NAND2X1 NAND2X1_1750 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf3_), .B(module_2_W_131_), .Y(_13036_) );
INVX1 INVX1_1884 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf2_), .Y(_13037_) );
NAND2X1 NAND2X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_13037_), .B(_12929_), .Y(_13038_) );
AOI21X1 AOI21X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_13038_), .B(_13036_), .C(module_2_W_179_), .Y(_13039_) );
INVX1 INVX1_1885 ( .gnd(gnd), .vdd(vdd), .A(_13039_), .Y(module_2_W_203_) );
XNOR2X1 XNOR2X1_354 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_132_), .B(bloque_datos_60_bF_buf1_), .Y(_13040_) );
NAND2X1 NAND2X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_13040_), .B(_12993_), .Y(module_2_W_204_) );
NAND2X1 NAND2X1_1753 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf3_), .B(module_2_W_133_), .Y(_13041_) );
OR2X2 OR2X2_311 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_133_), .B(bloque_datos_61_bF_buf2_), .Y(_13042_) );
AOI21X1 AOI21X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_13041_), .B(_13042_), .C(module_2_W_181_), .Y(_13043_) );
INVX1 INVX1_1886 ( .gnd(gnd), .vdd(vdd), .A(_13043_), .Y(module_2_W_205_) );
INVX2 INVX2_464 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf1_), .Y(_13044_) );
NAND2X1 NAND2X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_13044_), .B(_13001_), .Y(module_2_W_206_) );
INVX2 INVX2_465 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[63]), .Y(_13045_) );
NAND2X1 NAND2X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_13045_), .B(_13003_), .Y(module_2_W_207_) );
OAI21X1 OAI21X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_12943_), .B(bloque_datos_80_bF_buf1_), .C(bloque_datos_64_bF_buf3_), .Y(_13046_) );
OR2X2 OR2X2_312 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_136_), .B(bloque_datos_64_bF_buf2_), .Y(_13047_) );
AOI21X1 AOI21X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_13046_), .B(_13047_), .C(module_2_W_184_), .Y(_13048_) );
INVX1 INVX1_1887 ( .gnd(gnd), .vdd(vdd), .A(_13048_), .Y(module_2_W_208_) );
NAND2X1 NAND2X1_1756 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_65_bF_buf2_), .B(module_2_W_137_), .Y(_13049_) );
OR2X2 OR2X2_313 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_137_), .B(bloque_datos_65_bF_buf1_), .Y(_13050_) );
AOI21X1 AOI21X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_13049_), .B(_13050_), .C(module_2_W_185_), .Y(_13051_) );
INVX1 INVX1_1888 ( .gnd(gnd), .vdd(vdd), .A(_13051_), .Y(module_2_W_209_) );
OAI21X1 OAI21X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_12951_), .B(bloque_datos_82_bF_buf0_), .C(bloque_datos_66_bF_buf3_), .Y(_13052_) );
OR2X2 OR2X2_314 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_138_), .B(bloque_datos_66_bF_buf2_), .Y(_13053_) );
AOI21X1 AOI21X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_13052_), .B(_13053_), .C(module_2_W_186_), .Y(_13054_) );
INVX1 INVX1_1889 ( .gnd(gnd), .vdd(vdd), .A(_13054_), .Y(module_2_W_210_) );
OAI21X1 OAI21X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_12954_), .B(bloque_datos_83_bF_buf1_), .C(bloque_datos_67_bF_buf0_), .Y(_13055_) );
OR2X2 OR2X2_315 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_139_), .B(bloque_datos_67_bF_buf4_), .Y(_13056_) );
AOI21X1 AOI21X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_13055_), .B(_13056_), .C(module_2_W_187_), .Y(_13057_) );
INVX1 INVX1_1890 ( .gnd(gnd), .vdd(vdd), .A(_13057_), .Y(module_2_W_211_) );
NAND2X1 NAND2X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_12973_), .B(_13009_), .Y(module_2_W_212_) );
NAND2X1 NAND2X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_12976_), .B(_13011_), .Y(module_2_W_213_) );
NAND2X1 NAND2X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_12979_), .B(_13013_), .Y(module_2_W_214_) );
INVX1 INVX1_1891 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf0_), .Y(_13058_) );
NAND2X1 NAND2X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_13058_), .B(_13015_), .Y(module_2_W_215_) );
OR2X2 OR2X2_316 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_192_), .B(bloque_datos_72_bF_buf2_), .Y(module_2_W_216_) );
OR2X2 OR2X2_317 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_193_), .B(bloque_datos_73_bF_buf0_), .Y(module_2_W_217_) );
OR2X2 OR2X2_318 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_194_), .B(bloque_datos_74_bF_buf2_), .Y(module_2_W_218_) );
OR2X2 OR2X2_319 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_195_), .B(bloque_datos_75_bF_buf4_), .Y(module_2_W_219_) );
NAND2X1 NAND2X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_12932_), .B(_13022_), .Y(module_2_W_220_) );
NAND2X1 NAND2X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_12995_), .B(_13023_), .Y(module_2_W_221_) );
OR2X2 OR2X2_320 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_198_), .B(bloque_datos_78_bF_buf2_), .Y(module_2_W_222_) );
OR2X2 OR2X2_321 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_199_), .B(bloque_datos_79_bF_buf0_), .Y(module_2_W_223_) );
XNOR2X1 XNOR2X1_355 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_152_), .B(bloque_datos_80_bF_buf0_), .Y(_13059_) );
NAND2X1 NAND2X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_13028_), .B(_13059_), .Y(module_2_W_224_) );
OAI21X1 OAI21X1_2092 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_129_), .B(_12925_), .C(bloque_datos_81_bF_buf2_), .Y(_13060_) );
NAND3X1 NAND3X1_2939 ( .gnd(gnd), .vdd(vdd), .A(_12947_), .B(_12988_), .C(_12987_), .Y(_13061_) );
NAND2X1 NAND2X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_13060_), .B(_13061_), .Y(_13062_) );
NAND2X1 NAND2X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_13062_), .B(_13031_), .Y(module_2_W_225_) );
XNOR2X1 XNOR2X1_356 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_154_), .B(bloque_datos_82_bF_buf4_), .Y(_13063_) );
NAND2X1 NAND2X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_13035_), .B(_13063_), .Y(module_2_W_226_) );
XNOR2X1 XNOR2X1_357 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_155_), .B(bloque_datos_83_bF_buf0_), .Y(_13064_) );
NAND2X1 NAND2X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_13039_), .B(_13064_), .Y(module_2_W_227_) );
INVX1 INVX1_1892 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf2_), .Y(_13065_) );
NAND3X1 NAND3X1_2940 ( .gnd(gnd), .vdd(vdd), .A(_13065_), .B(_13040_), .C(_12993_), .Y(module_2_W_228_) );
OAI21X1 OAI21X1_2093 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_133_), .B(_12937_), .C(bloque_datos_85_bF_buf0_), .Y(_13066_) );
INVX1 INVX1_1893 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf4_), .Y(_13067_) );
NAND3X1 NAND3X1_2941 ( .gnd(gnd), .vdd(vdd), .A(_13067_), .B(_12998_), .C(_12997_), .Y(_13068_) );
NAND2X1 NAND2X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_13066_), .B(_13068_), .Y(_13069_) );
NAND2X1 NAND2X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_13069_), .B(_13043_), .Y(module_2_W_229_) );
INVX1 INVX1_1894 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf2_), .Y(_13070_) );
NAND3X1 NAND3X1_2942 ( .gnd(gnd), .vdd(vdd), .A(_13070_), .B(_13044_), .C(_13001_), .Y(module_2_W_230_) );
INVX1 INVX1_1895 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf1_), .Y(_13071_) );
NAND3X1 NAND3X1_2943 ( .gnd(gnd), .vdd(vdd), .A(_13071_), .B(_13045_), .C(_13003_), .Y(module_2_W_231_) );
AOI21X1 AOI21X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_12945_), .B(_12944_), .C(_12892_), .Y(_13072_) );
NOR2X1 NOR2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf4_), .B(module_2_W_160_), .Y(_13073_) );
OAI21X1 OAI21X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_13073_), .B(_13072_), .C(_13048_), .Y(module_2_W_232_) );
AOI21X1 AOI21X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_12950_), .B(_12949_), .C(_12896_), .Y(_13074_) );
NOR2X1 NOR2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf1_), .B(module_2_W_161_), .Y(_13075_) );
OAI21X1 OAI21X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_13074_), .B(_13075_), .C(_13051_), .Y(module_2_W_233_) );
AOI21X1 AOI21X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_12953_), .B(_12952_), .C(_12900_), .Y(_13076_) );
NOR2X1 NOR2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf4_), .B(module_2_W_162_), .Y(_13077_) );
OAI21X1 OAI21X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_13077_), .B(_13076_), .C(_13054_), .Y(module_2_W_234_) );
AOI21X1 AOI21X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_12956_), .B(_12955_), .C(_12904_), .Y(_13078_) );
NOR2X1 NOR2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf1_), .B(module_2_W_163_), .Y(_13079_) );
OAI21X1 OAI21X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_13079_), .B(_13078_), .C(_13057_), .Y(module_2_W_235_) );
NAND3X1 NAND3X1_2944 ( .gnd(gnd), .vdd(vdd), .A(_12908_), .B(_12973_), .C(_13009_), .Y(module_2_W_236_) );
NAND3X1 NAND3X1_2945 ( .gnd(gnd), .vdd(vdd), .A(_12912_), .B(_12976_), .C(_13011_), .Y(module_2_W_237_) );
NAND3X1 NAND3X1_2946 ( .gnd(gnd), .vdd(vdd), .A(_12916_), .B(_12979_), .C(_13013_), .Y(module_2_W_238_) );
NAND3X1 NAND3X1_2947 ( .gnd(gnd), .vdd(vdd), .A(_12920_), .B(_13058_), .C(_13015_), .Y(module_2_W_239_) );
OR2X2 OR2X2_322 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_192_), .B(module_2_W_128_), .Y(module_2_W_240_) );
OR2X2 OR2X2_323 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_193_), .B(module_2_W_129_), .Y(module_2_W_241_) );
OR2X2 OR2X2_324 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_194_), .B(module_2_W_130_), .Y(module_2_W_242_) );
OR2X2 OR2X2_325 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_195_), .B(module_2_W_131_), .Y(module_2_W_243_) );
NAND2X1 NAND2X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_12934_), .B(_13022_), .Y(module_2_W_244_) );
NAND2X1 NAND2X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_12997_), .B(_13023_), .Y(module_2_W_245_) );
OR2X2 OR2X2_326 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_198_), .B(module_2_W_134_), .Y(module_2_W_246_) );
OR2X2 OR2X2_327 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_199_), .B(module_2_W_135_), .Y(module_2_W_247_) );
XNOR2X1 XNOR2X1_358 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_176_), .B(module_2_W_136_), .Y(_13080_) );
NAND3X1 NAND3X1_2948 ( .gnd(gnd), .vdd(vdd), .A(_13028_), .B(_13059_), .C(_13080_), .Y(module_2_W_248_) );
NAND3X1 NAND3X1_2949 ( .gnd(gnd), .vdd(vdd), .A(_12949_), .B(_13062_), .C(_13031_), .Y(module_2_W_249_) );
XNOR2X1 XNOR2X1_359 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_178_), .B(module_2_W_138_), .Y(_13081_) );
NAND3X1 NAND3X1_2950 ( .gnd(gnd), .vdd(vdd), .A(_13035_), .B(_13063_), .C(_13081_), .Y(module_2_W_250_) );
XNOR2X1 XNOR2X1_360 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_179_), .B(module_2_W_139_), .Y(_13082_) );
NAND3X1 NAND3X1_2951 ( .gnd(gnd), .vdd(vdd), .A(_13039_), .B(_13064_), .C(_13082_), .Y(module_2_W_251_) );
INVX1 INVX1_1896 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_140_), .Y(_13083_) );
NAND3X1 NAND3X1_2952 ( .gnd(gnd), .vdd(vdd), .A(_13083_), .B(_13040_), .C(_12993_), .Y(module_2_W_252_) );
INVX1 INVX1_1897 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_141_), .Y(_13084_) );
NAND3X1 NAND3X1_2953 ( .gnd(gnd), .vdd(vdd), .A(_13084_), .B(_13069_), .C(_13043_), .Y(module_2_W_253_) );
INVX1 INVX1_1898 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_142_), .Y(_13085_) );
NAND3X1 NAND3X1_2954 ( .gnd(gnd), .vdd(vdd), .A(_13044_), .B(_13085_), .C(_13001_), .Y(module_2_W_254_) );
INVX1 INVX1_1899 ( .gnd(gnd), .vdd(vdd), .A(module_2_W_143_), .Y(_13086_) );
NAND3X1 NAND3X1_2955 ( .gnd(gnd), .vdd(vdd), .A(_13045_), .B(_13086_), .C(_13003_), .Y(module_2_W_255_) );
NAND3X1 NAND3X1_2956 ( .gnd(gnd), .vdd(vdd), .A(_13319_), .B(_13320_), .C(_13321_), .Y(_13322_) );
NAND2X1 NAND2X1_1772 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_200_), .B(_13304_), .Y(_13323_) );
OR2X2 OR2X2_328 ( .gnd(gnd), .vdd(vdd), .A(_13304_), .B(module_3_W_200_), .Y(_13324_) );
NAND2X1 NAND2X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_13323_), .B(_13324_), .Y(_13325_) );
NAND3X1 NAND3X1_2957 ( .gnd(gnd), .vdd(vdd), .A(_13322_), .B(_13325_), .C(_13317_), .Y(_13326_) );
NAND2X1 NAND2X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_13322_), .B(_13317_), .Y(_13327_) );
INVX2 INVX2_466 ( .gnd(gnd), .vdd(vdd), .A(_13325_), .Y(_13328_) );
AOI21X1 AOI21X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_13328_), .B(_13327_), .C(_15310_), .Y(_13329_) );
NAND3X1 NAND3X1_2958 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_228_), .B(_13326_), .C(_13329_), .Y(_13330_) );
INVX1 INVX1_1900 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_228_), .Y(_13331_) );
AOI21X1 AOI21X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_13320_), .B(_13321_), .C(_13319_), .Y(_13332_) );
NAND3X1 NAND3X1_2959 ( .gnd(gnd), .vdd(vdd), .A(_16739_), .B(_13312_), .C(_13309_), .Y(_13333_) );
NAND3X1 NAND3X1_2960 ( .gnd(gnd), .vdd(vdd), .A(_16742_), .B(_13314_), .C(_13315_), .Y(_13334_) );
AOI21X1 AOI21X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_13333_), .B(_13334_), .C(_16795_), .Y(_13335_) );
OAI21X1 OAI21X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_13332_), .B(_13335_), .C(_13328_), .Y(_13336_) );
NAND3X1 NAND3X1_2961 ( .gnd(gnd), .vdd(vdd), .A(_15299_), .B(_13326_), .C(_13336_), .Y(_13337_) );
NAND2X1 NAND2X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_13331_), .B(_13337_), .Y(_13338_) );
AOI21X1 AOI21X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_13338_), .B(_13330_), .C(_16751_), .Y(_13339_) );
INVX1 INVX1_1901 ( .gnd(gnd), .vdd(vdd), .A(_16751_), .Y(_13340_) );
NAND2X1 NAND2X1_1776 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_228_), .B(_13337_), .Y(_13341_) );
NAND3X1 NAND3X1_2962 ( .gnd(gnd), .vdd(vdd), .A(_13331_), .B(_13326_), .C(_13329_), .Y(_13342_) );
AOI21X1 AOI21X1_1877 ( .gnd(gnd), .vdd(vdd), .A(_13341_), .B(_13342_), .C(_13340_), .Y(_13343_) );
OAI21X1 OAI21X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_13339_), .B(_13343_), .C(_16793_), .Y(_13344_) );
OAI21X1 OAI21X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_16757_), .B(_16759_), .C(_16752_), .Y(_13345_) );
NAND3X1 NAND3X1_2963 ( .gnd(gnd), .vdd(vdd), .A(_13340_), .B(_13341_), .C(_13342_), .Y(_13346_) );
NAND3X1 NAND3X1_2964 ( .gnd(gnd), .vdd(vdd), .A(_16751_), .B(_13338_), .C(_13330_), .Y(_13347_) );
NAND3X1 NAND3X1_2965 ( .gnd(gnd), .vdd(vdd), .A(_13345_), .B(_13346_), .C(_13347_), .Y(_13348_) );
NAND2X1 NAND2X1_1777 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_216_), .B(_13325_), .Y(_13349_) );
OR2X2 OR2X2_329 ( .gnd(gnd), .vdd(vdd), .A(_13325_), .B(module_3_W_216_), .Y(_13350_) );
NAND2X1 NAND2X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_13349_), .B(_13350_), .Y(_13351_) );
NAND3X1 NAND3X1_2966 ( .gnd(gnd), .vdd(vdd), .A(_13348_), .B(_13351_), .C(_13344_), .Y(_13352_) );
AOI21X1 AOI21X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_13346_), .B(_13347_), .C(_13345_), .Y(_13353_) );
NOR3X1 NOR3X1_400 ( .gnd(gnd), .vdd(vdd), .A(_13339_), .B(_13343_), .C(_16793_), .Y(_13354_) );
INVX2 INVX2_467 ( .gnd(gnd), .vdd(vdd), .A(_13351_), .Y(_13355_) );
OAI21X1 OAI21X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_13354_), .B(_13353_), .C(_13355_), .Y(_13356_) );
NAND3X1 NAND3X1_2967 ( .gnd(gnd), .vdd(vdd), .A(_16544_), .B(_13352_), .C(_13356_), .Y(_13357_) );
NAND2X1 NAND2X1_1779 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_244_), .B(_13357_), .Y(_13358_) );
INVX1 INVX1_1902 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_244_), .Y(_13359_) );
NAND2X1 NAND2X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_13348_), .B(_13344_), .Y(_13360_) );
AOI21X1 AOI21X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_13355_), .B(_13360_), .C(_16545_), .Y(_13361_) );
NAND3X1 NAND3X1_2968 ( .gnd(gnd), .vdd(vdd), .A(_13359_), .B(_13352_), .C(_13361_), .Y(_13362_) );
NAND3X1 NAND3X1_2969 ( .gnd(gnd), .vdd(vdd), .A(_16792_), .B(_13362_), .C(_13358_), .Y(_13363_) );
NAND3X1 NAND3X1_2970 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_244_), .B(_13352_), .C(_13361_), .Y(_13364_) );
NAND2X1 NAND2X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_13359_), .B(_13357_), .Y(_13365_) );
NAND3X1 NAND3X1_2971 ( .gnd(gnd), .vdd(vdd), .A(_16764_), .B(_13364_), .C(_13365_), .Y(_13366_) );
AOI21X1 AOI21X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_13363_), .B(_13366_), .C(_16791_), .Y(_13367_) );
NOR2X1 NOR2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_16540_), .B(_16765_), .Y(_13368_) );
AOI21X1 AOI21X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_16555_), .B(_16768_), .C(_13368_), .Y(_13369_) );
AOI21X1 AOI21X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_13364_), .B(_13365_), .C(_16764_), .Y(_13370_) );
AOI21X1 AOI21X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_13362_), .B(_13358_), .C(_16792_), .Y(_13371_) );
NOR3X1 NOR3X1_401 ( .gnd(gnd), .vdd(vdd), .A(_13370_), .B(_13369_), .C(_13371_), .Y(_13372_) );
NOR2X1 NOR2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_232_), .B(_13355_), .Y(_13373_) );
AND2X2 AND2X2_304 ( .gnd(gnd), .vdd(vdd), .A(_13355_), .B(module_3_W_232_), .Y(_13374_) );
NOR2X1 NOR2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_13373_), .B(_13374_), .Y(_13375_) );
OAI21X1 OAI21X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_13372_), .B(_13367_), .C(_13375_), .Y(_13376_) );
OAI21X1 OAI21X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_13370_), .B(_13371_), .C(_13369_), .Y(_13377_) );
NAND3X1 NAND3X1_2972 ( .gnd(gnd), .vdd(vdd), .A(_13363_), .B(_13366_), .C(_16791_), .Y(_13378_) );
INVX2 INVX2_468 ( .gnd(gnd), .vdd(vdd), .A(_13375_), .Y(_13379_) );
NAND3X1 NAND3X1_2973 ( .gnd(gnd), .vdd(vdd), .A(_13379_), .B(_13378_), .C(_13377_), .Y(_13380_) );
NAND2X1 NAND2X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_13380_), .B(_13376_), .Y(_13381_) );
XNOR2X1 XNOR2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_13381_), .B(_16788_), .Y(module_3_H_4_) );
NAND3X1 NAND3X1_2974 ( .gnd(gnd), .vdd(vdd), .A(_16788_), .B(_13380_), .C(_13376_), .Y(_13382_) );
NOR2X1 NOR2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_216_), .B(_13328_), .Y(_13383_) );
NOR2X1 NOR2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_200_), .B(_13305_), .Y(_13384_) );
NOR2X1 NOR2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_184_), .B(_13280_), .Y(_13385_) );
INVX1 INVX1_1903 ( .gnd(gnd), .vdd(vdd), .A(_13258_), .Y(_13386_) );
NOR2X1 NOR2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_168_), .B(_13386_), .Y(_13387_) );
NOR2X1 NOR2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_152_), .B(_13236_), .Y(_13388_) );
INVX1 INVX1_1904 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_153_), .Y(_13389_) );
NOR2X1 NOR2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_136_), .B(_13213_), .Y(_13390_) );
INVX1 INVX1_1905 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_137_), .Y(_13391_) );
INVX1 INVX1_1906 ( .gnd(gnd), .vdd(vdd), .A(_13183_), .Y(_13392_) );
NOR2X1 NOR2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf3_), .B(_13392_), .Y(_13393_) );
INVX1 INVX1_1907 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf0_), .Y(_13394_) );
INVX1 INVX1_1908 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_73_bF_buf3_), .Y(_13395_) );
NOR2X1 NOR2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf1_), .B(_13133_), .Y(_13396_) );
NOR2X1 NOR2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf1_), .B(_13108_), .Y(_13397_) );
NOR2X1 NOR2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf1_), .B(_16894_), .Y(_13398_) );
NOR2X1 NOR2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .B(_16869_), .Y(_13399_) );
INVX1 INVX1_1909 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_25_), .Y(_13400_) );
INVX2 INVX2_469 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_9_), .Y(_13401_) );
NOR2X1 NOR2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_13400_), .B(_13401_), .Y(_13402_) );
NOR2X1 NOR2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_25_), .B(module_3_W_9_), .Y(_13403_) );
NOR2X1 NOR2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_13403_), .B(_13402_), .Y(_13404_) );
NOR2X1 NOR2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_16867_), .B(_13404_), .Y(_13405_) );
AND2X2 AND2X2_305 ( .gnd(gnd), .vdd(vdd), .A(_13404_), .B(_16867_), .Y(_13406_) );
NOR2X1 NOR2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_13405_), .B(_13406_), .Y(_13407_) );
NOR2X1 NOR2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .B(_13407_), .Y(_13408_) );
INVX1 INVX1_1910 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .Y(_13409_) );
OR2X2 OR2X2_330 ( .gnd(gnd), .vdd(vdd), .A(_13406_), .B(_13405_), .Y(_13410_) );
NOR2X1 NOR2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_13409_), .B(_13410_), .Y(_13411_) );
OAI21X1 OAI21X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_13411_), .B(_13408_), .C(_13399_), .Y(_13412_) );
OR2X2 OR2X2_331 ( .gnd(gnd), .vdd(vdd), .A(_13411_), .B(_13408_), .Y(_13413_) );
OR2X2 OR2X2_332 ( .gnd(gnd), .vdd(vdd), .A(_13413_), .B(_13399_), .Y(_13414_) );
AND2X2 AND2X2_306 ( .gnd(gnd), .vdd(vdd), .A(_13414_), .B(_13412_), .Y(_13415_) );
NOR2X1 NOR2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf0_), .B(_13415_), .Y(_13416_) );
AND2X2 AND2X2_307 ( .gnd(gnd), .vdd(vdd), .A(_13415_), .B(bloque_datos_25_bF_buf3_), .Y(_13417_) );
OAI21X1 OAI21X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_13417_), .B(_13416_), .C(_13398_), .Y(_13418_) );
OR2X2 OR2X2_333 ( .gnd(gnd), .vdd(vdd), .A(_13417_), .B(_13416_), .Y(_13419_) );
OR2X2 OR2X2_334 ( .gnd(gnd), .vdd(vdd), .A(_13419_), .B(_13398_), .Y(_13420_) );
AND2X2 AND2X2_308 ( .gnd(gnd), .vdd(vdd), .A(_13420_), .B(_13418_), .Y(_13421_) );
NOR2X1 NOR2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf0_), .B(_13421_), .Y(_13422_) );
INVX1 INVX1_1911 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf3_), .Y(_13423_) );
NAND2X1 NAND2X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_13418_), .B(_13420_), .Y(_13424_) );
NOR2X1 NOR2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_13423_), .B(_13424_), .Y(_13425_) );
OAI21X1 OAI21X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_13422_), .B(_13425_), .C(_13397_), .Y(_13426_) );
OR2X2 OR2X2_335 ( .gnd(gnd), .vdd(vdd), .A(_13422_), .B(_13425_), .Y(_13427_) );
OR2X2 OR2X2_336 ( .gnd(gnd), .vdd(vdd), .A(_13427_), .B(_13397_), .Y(_13428_) );
AND2X2 AND2X2_309 ( .gnd(gnd), .vdd(vdd), .A(_13428_), .B(_13426_), .Y(_13429_) );
NOR2X1 NOR2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf0_), .B(_13429_), .Y(_13430_) );
INVX1 INVX1_1912 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf3_), .Y(_13431_) );
NAND2X1 NAND2X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_13426_), .B(_13428_), .Y(_13432_) );
NOR2X1 NOR2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_13431_), .B(_13432_), .Y(_13433_) );
OAI21X1 OAI21X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_13430_), .B(_13433_), .C(_13396_), .Y(_13434_) );
OR2X2 OR2X2_337 ( .gnd(gnd), .vdd(vdd), .A(_13430_), .B(_13433_), .Y(_13435_) );
OR2X2 OR2X2_338 ( .gnd(gnd), .vdd(vdd), .A(_13435_), .B(_13396_), .Y(_13436_) );
NAND2X1 NAND2X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_13434_), .B(_13436_), .Y(_13437_) );
NAND2X1 NAND2X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_13395_), .B(_13437_), .Y(_13438_) );
OR2X2 OR2X2_339 ( .gnd(gnd), .vdd(vdd), .A(_13437_), .B(_13395_), .Y(_13439_) );
NAND2X1 NAND2X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_13438_), .B(_13439_), .Y(_13440_) );
NAND2X1 NAND2X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_13180_), .B(_13440_), .Y(_13441_) );
OR2X2 OR2X2_340 ( .gnd(gnd), .vdd(vdd), .A(_13440_), .B(_13180_), .Y(_13442_) );
NAND2X1 NAND2X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_13441_), .B(_13442_), .Y(_13443_) );
NAND2X1 NAND2X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_13394_), .B(_13443_), .Y(_13444_) );
OR2X2 OR2X2_341 ( .gnd(gnd), .vdd(vdd), .A(_13443_), .B(_13394_), .Y(_13445_) );
NAND2X1 NAND2X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_13444_), .B(_13445_), .Y(_13446_) );
NAND2X1 NAND2X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_13393_), .B(_13446_), .Y(_13447_) );
NOR2X1 NOR2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_13393_), .B(_13446_), .Y(_13448_) );
INVX1 INVX1_1913 ( .gnd(gnd), .vdd(vdd), .A(_13448_), .Y(_13449_) );
NAND2X1 NAND2X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_13447_), .B(_13449_), .Y(_13450_) );
NAND2X1 NAND2X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_13391_), .B(_13450_), .Y(_13451_) );
INVX2 INVX2_470 ( .gnd(gnd), .vdd(vdd), .A(_13450_), .Y(_13452_) );
NAND2X1 NAND2X1_1795 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_137_), .B(_13452_), .Y(_13453_) );
NAND2X1 NAND2X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_13451_), .B(_13453_), .Y(_13454_) );
NAND2X1 NAND2X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_13390_), .B(_13454_), .Y(_13455_) );
NOR2X1 NOR2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_13390_), .B(_13454_), .Y(_13456_) );
INVX1 INVX1_1914 ( .gnd(gnd), .vdd(vdd), .A(_13456_), .Y(_13457_) );
NAND2X1 NAND2X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_13455_), .B(_13457_), .Y(_13458_) );
NAND2X1 NAND2X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_13389_), .B(_13458_), .Y(_13459_) );
NOR2X1 NOR2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_13389_), .B(_13458_), .Y(_13460_) );
INVX1 INVX1_1915 ( .gnd(gnd), .vdd(vdd), .A(_13460_), .Y(_13461_) );
NAND2X1 NAND2X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_13459_), .B(_13461_), .Y(_13462_) );
NAND2X1 NAND2X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_13388_), .B(_13462_), .Y(_13463_) );
NOR2X1 NOR2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_13388_), .B(_13462_), .Y(_13464_) );
INVX1 INVX1_1916 ( .gnd(gnd), .vdd(vdd), .A(_13464_), .Y(_13465_) );
NAND2X1 NAND2X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_13463_), .B(_13465_), .Y(_13466_) );
INVX2 INVX2_471 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .Y(_13467_) );
NOR2X1 NOR2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_169_), .B(_13467_), .Y(_13468_) );
NAND2X1 NAND2X1_1803 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_169_), .B(_13467_), .Y(_13469_) );
INVX2 INVX2_472 ( .gnd(gnd), .vdd(vdd), .A(_13469_), .Y(_13470_) );
OAI21X1 OAI21X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_13470_), .B(_13468_), .C(_13387_), .Y(_13471_) );
NOR2X1 NOR2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_13468_), .B(_13470_), .Y(_13472_) );
OAI21X1 OAI21X1_2109 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_168_), .B(_13386_), .C(_13472_), .Y(_13473_) );
NAND2X1 NAND2X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_13471_), .B(_13473_), .Y(_13474_) );
INVX2 INVX2_473 ( .gnd(gnd), .vdd(vdd), .A(_13474_), .Y(_13475_) );
NOR2X1 NOR2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_185_), .B(_13475_), .Y(_13476_) );
NAND2X1 NAND2X1_1805 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_185_), .B(_13475_), .Y(_13477_) );
INVX2 INVX2_474 ( .gnd(gnd), .vdd(vdd), .A(_13477_), .Y(_13478_) );
OAI21X1 OAI21X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_13478_), .B(_13476_), .C(_13385_), .Y(_13479_) );
NOR2X1 NOR2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_13476_), .B(_13478_), .Y(_13480_) );
OAI21X1 OAI21X1_2111 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_184_), .B(_13280_), .C(_13480_), .Y(_13481_) );
NAND2X1 NAND2X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_13479_), .B(_13481_), .Y(_13482_) );
INVX2 INVX2_475 ( .gnd(gnd), .vdd(vdd), .A(_13482_), .Y(_13483_) );
NOR2X1 NOR2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_201_), .B(_13483_), .Y(_13484_) );
NAND2X1 NAND2X1_1807 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_201_), .B(_13483_), .Y(_13485_) );
INVX2 INVX2_476 ( .gnd(gnd), .vdd(vdd), .A(_13485_), .Y(_13486_) );
OAI21X1 OAI21X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_13486_), .B(_13484_), .C(_13384_), .Y(_13487_) );
NOR2X1 NOR2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_13484_), .B(_13486_), .Y(_13488_) );
OAI21X1 OAI21X1_2113 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_200_), .B(_13305_), .C(_13488_), .Y(_13489_) );
NAND2X1 NAND2X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_13487_), .B(_13489_), .Y(_13490_) );
INVX2 INVX2_477 ( .gnd(gnd), .vdd(vdd), .A(_13490_), .Y(_13491_) );
NOR2X1 NOR2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_217_), .B(_13491_), .Y(_13492_) );
NAND2X1 NAND2X1_1809 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_217_), .B(_13491_), .Y(_13493_) );
INVX2 INVX2_478 ( .gnd(gnd), .vdd(vdd), .A(_13493_), .Y(_13494_) );
OAI21X1 OAI21X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_13494_), .B(_13492_), .C(_13383_), .Y(_13495_) );
NOR2X1 NOR2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_13492_), .B(_13494_), .Y(_13496_) );
OAI21X1 OAI21X1_2115 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_216_), .B(_13328_), .C(_13496_), .Y(_13497_) );
NAND2X1 NAND2X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_13495_), .B(_13497_), .Y(_13498_) );
INVX2 INVX2_479 ( .gnd(gnd), .vdd(vdd), .A(_13498_), .Y(_13499_) );
NOR2X1 NOR2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_233_), .B(_13499_), .Y(_13500_) );
NAND2X1 NAND2X1_1811 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_233_), .B(_13499_), .Y(_13501_) );
INVX2 INVX2_480 ( .gnd(gnd), .vdd(vdd), .A(_13501_), .Y(_13502_) );
OAI21X1 OAI21X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_13502_), .B(_13500_), .C(_13373_), .Y(_13503_) );
NOR2X1 NOR2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_13500_), .B(_13502_), .Y(_13504_) );
OAI21X1 OAI21X1_2117 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_232_), .B(_13355_), .C(_13504_), .Y(_13505_) );
NAND2X1 NAND2X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_13503_), .B(_13505_), .Y(_13506_) );
OAI21X1 OAI21X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_13371_), .B(_13369_), .C(_13363_), .Y(_13507_) );
INVX1 INVX1_1917 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_245_), .Y(_13508_) );
AOI21X1 AOI21X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_13345_), .B(_13347_), .C(_13339_), .Y(_13509_) );
INVX2 INVX2_481 ( .gnd(gnd), .vdd(vdd), .A(_13341_), .Y(_13510_) );
INVX1 INVX1_1918 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_229_), .Y(_13511_) );
AOI21X1 AOI21X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_13319_), .B(_13321_), .C(_13313_), .Y(_13512_) );
INVX2 INVX2_482 ( .gnd(gnd), .vdd(vdd), .A(_13314_), .Y(_13513_) );
INVX1 INVX1_1919 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_213_), .Y(_13514_) );
AOI21X1 AOI21X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_13299_), .B(_13297_), .C(_13289_), .Y(_13515_) );
INVX2 INVX2_483 ( .gnd(gnd), .vdd(vdd), .A(_13293_), .Y(_13516_) );
INVX1 INVX1_1920 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_197_), .Y(_13517_) );
AOI21X1 AOI21X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_13273_), .B(_13271_), .C(_13266_), .Y(_13518_) );
INVX2 INVX2_484 ( .gnd(gnd), .vdd(vdd), .A(_13267_), .Y(_13519_) );
INVX1 INVX1_1921 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_181_), .Y(_13520_) );
AOI21X1 AOI21X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_16801_), .B(_13254_), .C(_13247_), .Y(_13521_) );
INVX2 INVX2_485 ( .gnd(gnd), .vdd(vdd), .A(_13249_), .Y(_13522_) );
INVX1 INVX1_1922 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_165_), .Y(_13523_) );
INVX1 INVX1_1923 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .Y(_13524_) );
AOI21X1 AOI21X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_13227_), .B(_13229_), .C(_13222_), .Y(_13525_) );
INVX1 INVX1_1924 ( .gnd(gnd), .vdd(vdd), .A(_13223_), .Y(_13526_) );
INVX1 INVX1_1925 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_149_), .Y(_13527_) );
AOI21X1 AOI21X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_13199_), .B(_16804_), .C(_13209_), .Y(_13528_) );
AOI21X1 AOI21X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_13172_), .B(_13173_), .C(_16806_), .Y(_13529_) );
AOI21X1 AOI21X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_13176_), .B(_13178_), .C(_13529_), .Y(_13530_) );
NOR3X1 NOR3X1_402 ( .gnd(gnd), .vdd(vdd), .A(_13140_), .B(_16658_), .C(_13144_), .Y(_13531_) );
OAI21X1 OAI21X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_13531_), .B(_16808_), .C(_13153_), .Y(_13532_) );
AOI21X1 AOI21X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_13122_), .B(_13123_), .C(_16812_), .Y(_13533_) );
AOI21X1 AOI21X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_13128_), .B(_13126_), .C(_13533_), .Y(_13534_) );
AOI21X1 AOI21X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_13097_), .B(_13098_), .C(_16816_), .Y(_13535_) );
AOI21X1 AOI21X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_13103_), .B(_13101_), .C(_13535_), .Y(_13536_) );
INVX1 INVX1_1926 ( .gnd(gnd), .vdd(vdd), .A(_16887_), .Y(_13537_) );
AOI21X1 AOI21X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_16886_), .B(_16888_), .C(_13537_), .Y(_13538_) );
INVX1 INVX1_1927 ( .gnd(gnd), .vdd(vdd), .A(_16863_), .Y(_13539_) );
AOI21X1 AOI21X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_16864_), .B(_16862_), .C(_13539_), .Y(_13540_) );
AOI21X1 AOI21X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_16836_), .B(_16835_), .C(_16595_), .Y(_13541_) );
NOR2X1 NOR2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_13541_), .B(_16847_), .Y(_13542_) );
INVX1 INVX1_1928 ( .gnd(gnd), .vdd(vdd), .A(_16835_), .Y(_13543_) );
NOR2X1 NOR2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_15694_), .B(_15683_), .Y(_13544_) );
INVX2 INVX2_486 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_5_), .Y(_13545_) );
XNOR2X1 XNOR2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_16827_), .B(_13545_), .Y(_13546_) );
NAND2X1 NAND2X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_13544_), .B(_13546_), .Y(_13547_) );
INVX1 INVX1_1929 ( .gnd(gnd), .vdd(vdd), .A(_13544_), .Y(_13548_) );
NOR2X1 NOR2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_5_), .B(_16827_), .Y(_13549_) );
NOR2X1 NOR2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_13545_), .B(_16824_), .Y(_13550_) );
OAI21X1 OAI21X1_2120 ( .gnd(gnd), .vdd(vdd), .A(_13550_), .B(_13549_), .C(_13548_), .Y(_13551_) );
NAND3X1 NAND3X1_2975 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_21_), .B(_13547_), .C(_13551_), .Y(_13552_) );
INVX1 INVX1_1930 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_21_), .Y(_13553_) );
OAI21X1 OAI21X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_13550_), .B(_13549_), .C(_13544_), .Y(_13554_) );
OAI21X1 OAI21X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_15683_), .B(_15694_), .C(_13546_), .Y(_13555_) );
NAND3X1 NAND3X1_2976 ( .gnd(gnd), .vdd(vdd), .A(_13553_), .B(_13555_), .C(_13554_), .Y(_13556_) );
NAND3X1 NAND3X1_2977 ( .gnd(gnd), .vdd(vdd), .A(_13543_), .B(_13552_), .C(_13556_), .Y(_13557_) );
NAND3X1 NAND3X1_2978 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_21_), .B(_13555_), .C(_13554_), .Y(_13558_) );
NAND3X1 NAND3X1_2979 ( .gnd(gnd), .vdd(vdd), .A(_13553_), .B(_13547_), .C(_13551_), .Y(_13559_) );
NAND3X1 NAND3X1_2980 ( .gnd(gnd), .vdd(vdd), .A(_16835_), .B(_13559_), .C(_13558_), .Y(_13560_) );
AND2X2 AND2X2_310 ( .gnd(gnd), .vdd(vdd), .A(_13557_), .B(_13560_), .Y(_13561_) );
NAND2X1 NAND2X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_13561_), .B(_13542_), .Y(_13562_) );
NAND2X1 NAND2X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_13560_), .B(_13557_), .Y(_13563_) );
OAI21X1 OAI21X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_13541_), .B(_16847_), .C(_13563_), .Y(_13564_) );
XNOR2X1 XNOR2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_15770_), .B(module_3_W_9_), .Y(_13565_) );
NAND3X1 NAND3X1_2981 ( .gnd(gnd), .vdd(vdd), .A(_13565_), .B(_13564_), .C(_13562_), .Y(_13566_) );
NAND2X1 NAND2X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_16834_), .B(_16838_), .Y(_13567_) );
NOR2X1 NOR2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_13563_), .B(_13567_), .Y(_13568_) );
NOR2X1 NOR2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_13561_), .B(_13542_), .Y(_13569_) );
INVX1 INVX1_1931 ( .gnd(gnd), .vdd(vdd), .A(_13565_), .Y(_13570_) );
OAI21X1 OAI21X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_13569_), .B(_13568_), .C(_13570_), .Y(_13571_) );
NAND3X1 NAND3X1_2982 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf3_), .B(_13566_), .C(_13571_), .Y(_13572_) );
INVX1 INVX1_1932 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf2_), .Y(_13573_) );
NAND3X1 NAND3X1_2983 ( .gnd(gnd), .vdd(vdd), .A(_13570_), .B(_13564_), .C(_13562_), .Y(_13574_) );
OAI21X1 OAI21X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_13569_), .B(_13568_), .C(_13565_), .Y(_13575_) );
NAND3X1 NAND3X1_2984 ( .gnd(gnd), .vdd(vdd), .A(_13573_), .B(_13574_), .C(_13575_), .Y(_13576_) );
NAND3X1 NAND3X1_2985 ( .gnd(gnd), .vdd(vdd), .A(_16850_), .B(_13572_), .C(_13576_), .Y(_13577_) );
NAND3X1 NAND3X1_2986 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf1_), .B(_13574_), .C(_13575_), .Y(_13578_) );
NAND3X1 NAND3X1_2987 ( .gnd(gnd), .vdd(vdd), .A(_13573_), .B(_13566_), .C(_13571_), .Y(_13579_) );
NAND3X1 NAND3X1_2988 ( .gnd(gnd), .vdd(vdd), .A(_16856_), .B(_13578_), .C(_13579_), .Y(_13580_) );
NAND3X1 NAND3X1_2989 ( .gnd(gnd), .vdd(vdd), .A(_13540_), .B(_13577_), .C(_13580_), .Y(_13581_) );
NAND2X1 NAND2X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_16863_), .B(_16865_), .Y(_13582_) );
NAND3X1 NAND3X1_2990 ( .gnd(gnd), .vdd(vdd), .A(_16856_), .B(_13572_), .C(_13576_), .Y(_13583_) );
NAND3X1 NAND3X1_2991 ( .gnd(gnd), .vdd(vdd), .A(_16850_), .B(_13578_), .C(_13579_), .Y(_13584_) );
NAND3X1 NAND3X1_2992 ( .gnd(gnd), .vdd(vdd), .A(_13583_), .B(_13584_), .C(_13582_), .Y(_13585_) );
XNOR2X1 XNOR2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_15814_), .B(_13407_), .Y(_13586_) );
INVX1 INVX1_1933 ( .gnd(gnd), .vdd(vdd), .A(_13586_), .Y(_13587_) );
NAND3X1 NAND3X1_2993 ( .gnd(gnd), .vdd(vdd), .A(_13581_), .B(_13587_), .C(_13585_), .Y(_13588_) );
AOI21X1 AOI21X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_13583_), .B(_13584_), .C(_13582_), .Y(_13589_) );
AOI21X1 AOI21X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_13577_), .B(_13580_), .C(_13540_), .Y(_13590_) );
OAI21X1 OAI21X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_13589_), .B(_13590_), .C(_13586_), .Y(_13591_) );
NAND3X1 NAND3X1_2994 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf3_), .B(_13588_), .C(_13591_), .Y(_13592_) );
INVX1 INVX1_1934 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf2_), .Y(_13593_) );
NAND3X1 NAND3X1_2995 ( .gnd(gnd), .vdd(vdd), .A(_13581_), .B(_13586_), .C(_13585_), .Y(_13594_) );
OAI21X1 OAI21X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_13589_), .B(_13590_), .C(_13587_), .Y(_13595_) );
NAND3X1 NAND3X1_2996 ( .gnd(gnd), .vdd(vdd), .A(_13593_), .B(_13594_), .C(_13595_), .Y(_13596_) );
NAND3X1 NAND3X1_2997 ( .gnd(gnd), .vdd(vdd), .A(_16876_), .B(_13592_), .C(_13596_), .Y(_13597_) );
NAND3X1 NAND3X1_2998 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf1_), .B(_13594_), .C(_13595_), .Y(_13598_) );
NAND3X1 NAND3X1_2999 ( .gnd(gnd), .vdd(vdd), .A(_13593_), .B(_13588_), .C(_13591_), .Y(_13599_) );
NAND3X1 NAND3X1_3000 ( .gnd(gnd), .vdd(vdd), .A(_16882_), .B(_13598_), .C(_13599_), .Y(_13600_) );
NAND3X1 NAND3X1_3001 ( .gnd(gnd), .vdd(vdd), .A(_13597_), .B(_13600_), .C(_13538_), .Y(_13601_) );
INVX1 INVX1_1935 ( .gnd(gnd), .vdd(vdd), .A(_16888_), .Y(_13602_) );
OAI21X1 OAI21X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_13602_), .B(_16817_), .C(_16887_), .Y(_13603_) );
NAND3X1 NAND3X1_3002 ( .gnd(gnd), .vdd(vdd), .A(_16882_), .B(_13592_), .C(_13596_), .Y(_13604_) );
NAND3X1 NAND3X1_3003 ( .gnd(gnd), .vdd(vdd), .A(_16876_), .B(_13598_), .C(_13599_), .Y(_13605_) );
NAND3X1 NAND3X1_3004 ( .gnd(gnd), .vdd(vdd), .A(_13604_), .B(_13603_), .C(_13605_), .Y(_13606_) );
NAND2X1 NAND2X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_13412_), .B(_13414_), .Y(_13607_) );
XNOR2X1 XNOR2X1_365 ( .gnd(gnd), .vdd(vdd), .A(_15869_), .B(_13607_), .Y(_13608_) );
INVX1 INVX1_1936 ( .gnd(gnd), .vdd(vdd), .A(_13608_), .Y(_13609_) );
NAND3X1 NAND3X1_3005 ( .gnd(gnd), .vdd(vdd), .A(_13609_), .B(_13606_), .C(_13601_), .Y(_13610_) );
AOI21X1 AOI21X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_13604_), .B(_13605_), .C(_13603_), .Y(_13611_) );
AOI21X1 AOI21X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_13597_), .B(_13600_), .C(_13538_), .Y(_13612_) );
OAI21X1 OAI21X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_13611_), .B(_13612_), .C(_13608_), .Y(_13613_) );
NAND3X1 NAND3X1_3006 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf0_), .B(_13610_), .C(_13613_), .Y(_13614_) );
INVX1 INVX1_1937 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf3_), .Y(_13615_) );
NAND3X1 NAND3X1_3007 ( .gnd(gnd), .vdd(vdd), .A(_13608_), .B(_13606_), .C(_13601_), .Y(_13616_) );
OAI21X1 OAI21X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_13611_), .B(_13612_), .C(_13609_), .Y(_13617_) );
NAND3X1 NAND3X1_3008 ( .gnd(gnd), .vdd(vdd), .A(_13615_), .B(_13616_), .C(_13617_), .Y(_13618_) );
NAND3X1 NAND3X1_3009 ( .gnd(gnd), .vdd(vdd), .A(_13091_), .B(_13614_), .C(_13618_), .Y(_13619_) );
NAND3X1 NAND3X1_3010 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf2_), .B(_13616_), .C(_13617_), .Y(_13620_) );
NAND3X1 NAND3X1_3011 ( .gnd(gnd), .vdd(vdd), .A(_13615_), .B(_13610_), .C(_13613_), .Y(_13621_) );
NAND3X1 NAND3X1_3012 ( .gnd(gnd), .vdd(vdd), .A(_13097_), .B(_13620_), .C(_13621_), .Y(_13622_) );
NAND3X1 NAND3X1_3013 ( .gnd(gnd), .vdd(vdd), .A(_13536_), .B(_13619_), .C(_13622_), .Y(_13623_) );
NOR3X1 NOR3X1_403 ( .gnd(gnd), .vdd(vdd), .A(_13091_), .B(_16634_), .C(_13095_), .Y(_13624_) );
OAI21X1 OAI21X1_2131 ( .gnd(gnd), .vdd(vdd), .A(_13624_), .B(_16815_), .C(_13102_), .Y(_13625_) );
NAND3X1 NAND3X1_3014 ( .gnd(gnd), .vdd(vdd), .A(_13097_), .B(_13614_), .C(_13618_), .Y(_13626_) );
NAND3X1 NAND3X1_3015 ( .gnd(gnd), .vdd(vdd), .A(_13091_), .B(_13620_), .C(_13621_), .Y(_13627_) );
NAND3X1 NAND3X1_3016 ( .gnd(gnd), .vdd(vdd), .A(_13625_), .B(_13626_), .C(_13627_), .Y(_13628_) );
XNOR2X1 XNOR2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_15946_), .B(_13421_), .Y(_13629_) );
NAND3X1 NAND3X1_3017 ( .gnd(gnd), .vdd(vdd), .A(_13629_), .B(_13623_), .C(_13628_), .Y(_13630_) );
AOI21X1 AOI21X1_1904 ( .gnd(gnd), .vdd(vdd), .A(_13626_), .B(_13627_), .C(_13625_), .Y(_13631_) );
AOI21X1 AOI21X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_13619_), .B(_13622_), .C(_13536_), .Y(_13632_) );
INVX1 INVX1_1938 ( .gnd(gnd), .vdd(vdd), .A(_13629_), .Y(_13633_) );
OAI21X1 OAI21X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_13631_), .B(_13632_), .C(_13633_), .Y(_13634_) );
NAND3X1 NAND3X1_3018 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf0_), .B(_13630_), .C(_13634_), .Y(_13635_) );
INVX1 INVX1_1939 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf3_), .Y(_13636_) );
NAND3X1 NAND3X1_3019 ( .gnd(gnd), .vdd(vdd), .A(_13633_), .B(_13623_), .C(_13628_), .Y(_13637_) );
OAI21X1 OAI21X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_13631_), .B(_13632_), .C(_13629_), .Y(_13638_) );
NAND3X1 NAND3X1_3020 ( .gnd(gnd), .vdd(vdd), .A(_13636_), .B(_13637_), .C(_13638_), .Y(_13639_) );
NAND3X1 NAND3X1_3021 ( .gnd(gnd), .vdd(vdd), .A(_13115_), .B(_13635_), .C(_13639_), .Y(_13640_) );
NAND3X1 NAND3X1_3022 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf2_), .B(_13637_), .C(_13638_), .Y(_13641_) );
NAND3X1 NAND3X1_3023 ( .gnd(gnd), .vdd(vdd), .A(_13636_), .B(_13630_), .C(_13634_), .Y(_13642_) );
NAND3X1 NAND3X1_3024 ( .gnd(gnd), .vdd(vdd), .A(_13122_), .B(_13641_), .C(_13642_), .Y(_13643_) );
NAND3X1 NAND3X1_3025 ( .gnd(gnd), .vdd(vdd), .A(_13534_), .B(_13640_), .C(_13643_), .Y(_13644_) );
NOR3X1 NOR3X1_404 ( .gnd(gnd), .vdd(vdd), .A(_13115_), .B(_13121_), .C(_13119_), .Y(_13645_) );
OAI21X1 OAI21X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_13645_), .B(_16810_), .C(_13127_), .Y(_13646_) );
NAND3X1 NAND3X1_3026 ( .gnd(gnd), .vdd(vdd), .A(_13122_), .B(_13635_), .C(_13639_), .Y(_13647_) );
NAND3X1 NAND3X1_3027 ( .gnd(gnd), .vdd(vdd), .A(_13115_), .B(_13641_), .C(_13642_), .Y(_13648_) );
NAND3X1 NAND3X1_3028 ( .gnd(gnd), .vdd(vdd), .A(_13647_), .B(_13648_), .C(_13646_), .Y(_13649_) );
XNOR2X1 XNOR2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_16012_), .B(_13429_), .Y(_13650_) );
INVX1 INVX1_1940 ( .gnd(gnd), .vdd(vdd), .A(_13650_), .Y(_13651_) );
NAND3X1 NAND3X1_3029 ( .gnd(gnd), .vdd(vdd), .A(_13651_), .B(_13644_), .C(_13649_), .Y(_13652_) );
AOI21X1 AOI21X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_13647_), .B(_13648_), .C(_13646_), .Y(_13653_) );
AOI21X1 AOI21X1_1907 ( .gnd(gnd), .vdd(vdd), .A(_13640_), .B(_13643_), .C(_13534_), .Y(_13654_) );
OAI21X1 OAI21X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_13653_), .B(_13654_), .C(_13650_), .Y(_13655_) );
NAND3X1 NAND3X1_3030 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf0_), .B(_13652_), .C(_13655_), .Y(_13656_) );
INVX1 INVX1_1941 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf3_), .Y(_13657_) );
NAND3X1 NAND3X1_3031 ( .gnd(gnd), .vdd(vdd), .A(_13650_), .B(_13644_), .C(_13649_), .Y(_13658_) );
OAI21X1 OAI21X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_13653_), .B(_13654_), .C(_13651_), .Y(_13659_) );
NAND3X1 NAND3X1_3032 ( .gnd(gnd), .vdd(vdd), .A(_13657_), .B(_13658_), .C(_13659_), .Y(_13660_) );
NAND3X1 NAND3X1_3033 ( .gnd(gnd), .vdd(vdd), .A(_13146_), .B(_13656_), .C(_13660_), .Y(_13661_) );
NAND3X1 NAND3X1_3034 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf2_), .B(_13658_), .C(_13659_), .Y(_13662_) );
NAND3X1 NAND3X1_3035 ( .gnd(gnd), .vdd(vdd), .A(_13657_), .B(_13652_), .C(_13655_), .Y(_13663_) );
NAND3X1 NAND3X1_3036 ( .gnd(gnd), .vdd(vdd), .A(_13140_), .B(_13662_), .C(_13663_), .Y(_13664_) );
AOI21X1 AOI21X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_13661_), .B(_13664_), .C(_13532_), .Y(_13665_) );
AOI21X1 AOI21X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_13146_), .B(_13147_), .C(_16809_), .Y(_13666_) );
AOI21X1 AOI21X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_13152_), .B(_13154_), .C(_13666_), .Y(_13667_) );
NAND3X1 NAND3X1_3037 ( .gnd(gnd), .vdd(vdd), .A(_13140_), .B(_13656_), .C(_13660_), .Y(_13668_) );
NAND3X1 NAND3X1_3038 ( .gnd(gnd), .vdd(vdd), .A(_13146_), .B(_13662_), .C(_13663_), .Y(_13669_) );
AOI21X1 AOI21X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_13668_), .B(_13669_), .C(_13667_), .Y(_13670_) );
XNOR2X1 XNOR2X1_368 ( .gnd(gnd), .vdd(vdd), .A(_16056_), .B(_13437_), .Y(_13671_) );
NOR3X1 NOR3X1_405 ( .gnd(gnd), .vdd(vdd), .A(_13670_), .B(_13671_), .C(_13665_), .Y(_13672_) );
NAND3X1 NAND3X1_3039 ( .gnd(gnd), .vdd(vdd), .A(_13667_), .B(_13668_), .C(_13669_), .Y(_13673_) );
NAND3X1 NAND3X1_3040 ( .gnd(gnd), .vdd(vdd), .A(_13661_), .B(_13664_), .C(_13532_), .Y(_13674_) );
INVX1 INVX1_1942 ( .gnd(gnd), .vdd(vdd), .A(_13671_), .Y(_13675_) );
AOI21X1 AOI21X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_13673_), .B(_13674_), .C(_13675_), .Y(_13676_) );
OAI21X1 OAI21X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_13672_), .B(_13676_), .C(bloque_datos_85_bF_buf3_), .Y(_13677_) );
INVX1 INVX1_1943 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf2_), .Y(_13678_) );
NAND3X1 NAND3X1_3041 ( .gnd(gnd), .vdd(vdd), .A(_13675_), .B(_13673_), .C(_13674_), .Y(_13679_) );
OAI21X1 OAI21X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_13665_), .B(_13670_), .C(_13671_), .Y(_13680_) );
NAND3X1 NAND3X1_3042 ( .gnd(gnd), .vdd(vdd), .A(_13678_), .B(_13679_), .C(_13680_), .Y(_13681_) );
NAND3X1 NAND3X1_3043 ( .gnd(gnd), .vdd(vdd), .A(_13166_), .B(_13681_), .C(_13677_), .Y(_13682_) );
NAND3X1 NAND3X1_3044 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf1_), .B(_13679_), .C(_13680_), .Y(_13683_) );
OAI21X1 OAI21X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_13672_), .B(_13676_), .C(_13678_), .Y(_13684_) );
NAND3X1 NAND3X1_3045 ( .gnd(gnd), .vdd(vdd), .A(_13172_), .B(_13683_), .C(_13684_), .Y(_13685_) );
NAND3X1 NAND3X1_3046 ( .gnd(gnd), .vdd(vdd), .A(_13530_), .B(_13682_), .C(_13685_), .Y(_13686_) );
NOR3X1 NOR3X1_406 ( .gnd(gnd), .vdd(vdd), .A(_13166_), .B(_16670_), .C(_13170_), .Y(_13687_) );
OAI21X1 OAI21X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_13687_), .B(_16805_), .C(_13177_), .Y(_13688_) );
NAND3X1 NAND3X1_3047 ( .gnd(gnd), .vdd(vdd), .A(_13172_), .B(_13681_), .C(_13677_), .Y(_13689_) );
NAND3X1 NAND3X1_3048 ( .gnd(gnd), .vdd(vdd), .A(_13166_), .B(_13683_), .C(_13684_), .Y(_13690_) );
NAND3X1 NAND3X1_3049 ( .gnd(gnd), .vdd(vdd), .A(_13689_), .B(_13690_), .C(_13688_), .Y(_13691_) );
XNOR2X1 XNOR2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_16154_), .B(_13443_), .Y(_13692_) );
NAND3X1 NAND3X1_3050 ( .gnd(gnd), .vdd(vdd), .A(_13692_), .B(_13686_), .C(_13691_), .Y(_13693_) );
AOI21X1 AOI21X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_13689_), .B(_13690_), .C(_13688_), .Y(_13694_) );
AOI21X1 AOI21X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_13682_), .B(_13685_), .C(_13530_), .Y(_13695_) );
INVX1 INVX1_1944 ( .gnd(gnd), .vdd(vdd), .A(_13692_), .Y(_13696_) );
OAI21X1 OAI21X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_13694_), .B(_13695_), .C(_13696_), .Y(_13697_) );
NAND3X1 NAND3X1_3051 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_133_), .B(_13693_), .C(_13697_), .Y(_13698_) );
INVX1 INVX1_1945 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_133_), .Y(_13699_) );
NAND3X1 NAND3X1_3052 ( .gnd(gnd), .vdd(vdd), .A(_13696_), .B(_13686_), .C(_13691_), .Y(_13700_) );
OAI21X1 OAI21X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_13694_), .B(_13695_), .C(_13692_), .Y(_13701_) );
NAND3X1 NAND3X1_3053 ( .gnd(gnd), .vdd(vdd), .A(_13699_), .B(_13700_), .C(_13701_), .Y(_13702_) );
AOI21X1 AOI21X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_13698_), .B(_13702_), .C(_13190_), .Y(_13703_) );
NAND3X1 NAND3X1_3054 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_133_), .B(_13700_), .C(_13701_), .Y(_13704_) );
NAND3X1 NAND3X1_3055 ( .gnd(gnd), .vdd(vdd), .A(_13699_), .B(_13693_), .C(_13697_), .Y(_13705_) );
AOI21X1 AOI21X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_13704_), .B(_13705_), .C(_13197_), .Y(_13706_) );
OAI21X1 OAI21X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_13703_), .B(_13706_), .C(_13528_), .Y(_13707_) );
OAI21X1 OAI21X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_13210_), .B(_13201_), .C(_13195_), .Y(_13708_) );
AOI21X1 AOI21X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_13698_), .B(_13702_), .C(_13197_), .Y(_13709_) );
AOI21X1 AOI21X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_13704_), .B(_13705_), .C(_13190_), .Y(_13710_) );
OAI21X1 OAI21X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_13709_), .B(_13710_), .C(_13708_), .Y(_13711_) );
NAND3X1 NAND3X1_3056 ( .gnd(gnd), .vdd(vdd), .A(_13452_), .B(_13707_), .C(_13711_), .Y(_13712_) );
NAND3X1 NAND3X1_3057 ( .gnd(gnd), .vdd(vdd), .A(_13197_), .B(_13704_), .C(_13705_), .Y(_13713_) );
NAND3X1 NAND3X1_3058 ( .gnd(gnd), .vdd(vdd), .A(_13190_), .B(_13698_), .C(_13702_), .Y(_13714_) );
AOI21X1 AOI21X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_13713_), .B(_13714_), .C(_13708_), .Y(_13715_) );
NAND3X1 NAND3X1_3059 ( .gnd(gnd), .vdd(vdd), .A(_13190_), .B(_13704_), .C(_13705_), .Y(_13716_) );
NAND3X1 NAND3X1_3060 ( .gnd(gnd), .vdd(vdd), .A(_13197_), .B(_13698_), .C(_13702_), .Y(_13717_) );
AOI21X1 AOI21X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_13716_), .B(_13717_), .C(_13528_), .Y(_13718_) );
OAI21X1 OAI21X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_13715_), .B(_13718_), .C(_13450_), .Y(_13719_) );
NAND2X1 NAND2X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_13712_), .B(_13719_), .Y(_13720_) );
NAND3X1 NAND3X1_3061 ( .gnd(gnd), .vdd(vdd), .A(_13527_), .B(_16231_), .C(_13720_), .Y(_13721_) );
OAI21X1 OAI21X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_13715_), .B(_13718_), .C(_13452_), .Y(_13722_) );
NAND3X1 NAND3X1_3062 ( .gnd(gnd), .vdd(vdd), .A(_13450_), .B(_13707_), .C(_13711_), .Y(_13723_) );
NAND3X1 NAND3X1_3063 ( .gnd(gnd), .vdd(vdd), .A(_16231_), .B(_13723_), .C(_13722_), .Y(_13724_) );
NAND2X1 NAND2X1_1820 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_149_), .B(_13724_), .Y(_13725_) );
NAND3X1 NAND3X1_3064 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_13721_), .C(_13725_), .Y(_13726_) );
NOR2X1 NOR2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_149_), .B(_13724_), .Y(_13727_) );
AOI21X1 AOI21X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_16231_), .B(_13720_), .C(_13527_), .Y(_13728_) );
OAI21X1 OAI21X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_13727_), .B(_13728_), .C(_13223_), .Y(_13729_) );
NAND3X1 NAND3X1_3065 ( .gnd(gnd), .vdd(vdd), .A(_13726_), .B(_13525_), .C(_13729_), .Y(_13730_) );
OAI21X1 OAI21X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_13225_), .B(_16803_), .C(_13228_), .Y(_13731_) );
OAI21X1 OAI21X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_13727_), .B(_13728_), .C(_13526_), .Y(_13732_) );
NAND3X1 NAND3X1_3066 ( .gnd(gnd), .vdd(vdd), .A(_13223_), .B(_13721_), .C(_13725_), .Y(_13733_) );
NAND3X1 NAND3X1_3067 ( .gnd(gnd), .vdd(vdd), .A(_13733_), .B(_13732_), .C(_13731_), .Y(_13734_) );
NAND3X1 NAND3X1_3068 ( .gnd(gnd), .vdd(vdd), .A(_13524_), .B(_13730_), .C(_13734_), .Y(_13735_) );
AOI21X1 AOI21X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_13733_), .B(_13732_), .C(_13731_), .Y(_13736_) );
AOI21X1 AOI21X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_13726_), .B(_13729_), .C(_13525_), .Y(_13737_) );
OAI21X1 OAI21X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_13736_), .B(_13737_), .C(_13458_), .Y(_13738_) );
NAND2X1 NAND2X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_13735_), .B(_13738_), .Y(_13739_) );
NAND3X1 NAND3X1_3069 ( .gnd(gnd), .vdd(vdd), .A(_13523_), .B(_16315_), .C(_13739_), .Y(_13740_) );
OAI21X1 OAI21X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_13736_), .B(_13737_), .C(_13524_), .Y(_13741_) );
NAND3X1 NAND3X1_3070 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .B(_13730_), .C(_13734_), .Y(_13742_) );
NAND3X1 NAND3X1_3071 ( .gnd(gnd), .vdd(vdd), .A(_16315_), .B(_13742_), .C(_13741_), .Y(_13743_) );
NAND2X1 NAND2X1_1822 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_165_), .B(_13743_), .Y(_13744_) );
NAND3X1 NAND3X1_3072 ( .gnd(gnd), .vdd(vdd), .A(_13522_), .B(_13740_), .C(_13744_), .Y(_13745_) );
NOR2X1 NOR2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_165_), .B(_13743_), .Y(_13746_) );
AOI21X1 AOI21X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_16315_), .B(_13739_), .C(_13523_), .Y(_13747_) );
OAI21X1 OAI21X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_13746_), .B(_13747_), .C(_13249_), .Y(_13748_) );
NAND3X1 NAND3X1_3073 ( .gnd(gnd), .vdd(vdd), .A(_13521_), .B(_13745_), .C(_13748_), .Y(_13749_) );
OAI21X1 OAI21X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_16802_), .B(_13251_), .C(_13253_), .Y(_13750_) );
OAI21X1 OAI21X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_13746_), .B(_13747_), .C(_13522_), .Y(_13751_) );
NAND3X1 NAND3X1_3074 ( .gnd(gnd), .vdd(vdd), .A(_13249_), .B(_13740_), .C(_13744_), .Y(_13752_) );
NAND3X1 NAND3X1_3075 ( .gnd(gnd), .vdd(vdd), .A(_13752_), .B(_13750_), .C(_13751_), .Y(_13753_) );
NAND3X1 NAND3X1_3076 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .B(_13749_), .C(_13753_), .Y(_13754_) );
NAND2X1 NAND2X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_13749_), .B(_13753_), .Y(_13755_) );
AOI21X1 AOI21X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_13467_), .B(_13755_), .C(_16324_), .Y(_13756_) );
NAND3X1 NAND3X1_3077 ( .gnd(gnd), .vdd(vdd), .A(_13520_), .B(_13754_), .C(_13756_), .Y(_13757_) );
AOI21X1 AOI21X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_13752_), .B(_13751_), .C(_13750_), .Y(_13758_) );
AOI21X1 AOI21X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_13745_), .B(_13748_), .C(_13521_), .Y(_13759_) );
OAI21X1 OAI21X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_13758_), .B(_13759_), .C(_13467_), .Y(_13760_) );
NAND3X1 NAND3X1_3078 ( .gnd(gnd), .vdd(vdd), .A(_16323_), .B(_13754_), .C(_13760_), .Y(_13761_) );
NAND2X1 NAND2X1_1824 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_181_), .B(_13761_), .Y(_13762_) );
NAND3X1 NAND3X1_3079 ( .gnd(gnd), .vdd(vdd), .A(_13519_), .B(_13757_), .C(_13762_), .Y(_13763_) );
NOR2X1 NOR2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_181_), .B(_13761_), .Y(_13764_) );
AOI21X1 AOI21X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_13754_), .B(_13756_), .C(_13520_), .Y(_13765_) );
OAI21X1 OAI21X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_13764_), .B(_13765_), .C(_13267_), .Y(_13766_) );
NAND3X1 NAND3X1_3080 ( .gnd(gnd), .vdd(vdd), .A(_13518_), .B(_13763_), .C(_13766_), .Y(_13767_) );
OAI21X1 OAI21X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_13269_), .B(_16799_), .C(_13272_), .Y(_13768_) );
OAI21X1 OAI21X1_2159 ( .gnd(gnd), .vdd(vdd), .A(_13764_), .B(_13765_), .C(_13519_), .Y(_13769_) );
NAND3X1 NAND3X1_3081 ( .gnd(gnd), .vdd(vdd), .A(_13267_), .B(_13757_), .C(_13762_), .Y(_13770_) );
NAND3X1 NAND3X1_3082 ( .gnd(gnd), .vdd(vdd), .A(_13770_), .B(_13768_), .C(_13769_), .Y(_13771_) );
NAND3X1 NAND3X1_3083 ( .gnd(gnd), .vdd(vdd), .A(_13475_), .B(_13767_), .C(_13771_), .Y(_13772_) );
AOI21X1 AOI21X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_13770_), .B(_13769_), .C(_13768_), .Y(_13773_) );
AOI21X1 AOI21X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_13763_), .B(_13766_), .C(_13518_), .Y(_13774_) );
OAI21X1 OAI21X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_13773_), .B(_13774_), .C(_13474_), .Y(_13775_) );
NAND2X1 NAND2X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_13772_), .B(_13775_), .Y(_13776_) );
NAND3X1 NAND3X1_3084 ( .gnd(gnd), .vdd(vdd), .A(_13517_), .B(_16332_), .C(_13776_), .Y(_13777_) );
OAI21X1 OAI21X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_13773_), .B(_13774_), .C(_13475_), .Y(_13778_) );
NAND3X1 NAND3X1_3085 ( .gnd(gnd), .vdd(vdd), .A(_13474_), .B(_13767_), .C(_13771_), .Y(_13779_) );
NAND3X1 NAND3X1_3086 ( .gnd(gnd), .vdd(vdd), .A(_16332_), .B(_13779_), .C(_13778_), .Y(_13780_) );
NAND2X1 NAND2X1_1826 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_197_), .B(_13780_), .Y(_13781_) );
NAND3X1 NAND3X1_3087 ( .gnd(gnd), .vdd(vdd), .A(_13516_), .B(_13777_), .C(_13781_), .Y(_13782_) );
NOR2X1 NOR2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_197_), .B(_13780_), .Y(_13783_) );
AOI21X1 AOI21X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_16332_), .B(_13776_), .C(_13517_), .Y(_13784_) );
OAI21X1 OAI21X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_13783_), .B(_13784_), .C(_13293_), .Y(_13785_) );
NAND3X1 NAND3X1_3088 ( .gnd(gnd), .vdd(vdd), .A(_13782_), .B(_13515_), .C(_13785_), .Y(_13786_) );
OAI21X1 OAI21X1_2163 ( .gnd(gnd), .vdd(vdd), .A(_13295_), .B(_16797_), .C(_13298_), .Y(_13787_) );
OAI21X1 OAI21X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_13783_), .B(_13784_), .C(_13516_), .Y(_13788_) );
NAND3X1 NAND3X1_3089 ( .gnd(gnd), .vdd(vdd), .A(_13293_), .B(_13777_), .C(_13781_), .Y(_13789_) );
NAND3X1 NAND3X1_3090 ( .gnd(gnd), .vdd(vdd), .A(_13789_), .B(_13788_), .C(_13787_), .Y(_13790_) );
NAND3X1 NAND3X1_3091 ( .gnd(gnd), .vdd(vdd), .A(_13483_), .B(_13786_), .C(_13790_), .Y(_13791_) );
AOI21X1 AOI21X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_13789_), .B(_13788_), .C(_13787_), .Y(_13792_) );
AOI21X1 AOI21X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_13782_), .B(_13785_), .C(_13515_), .Y(_13793_) );
OAI21X1 OAI21X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_13792_), .B(_13793_), .C(_13482_), .Y(_13794_) );
NAND2X1 NAND2X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_13791_), .B(_13794_), .Y(_13795_) );
NAND3X1 NAND3X1_3092 ( .gnd(gnd), .vdd(vdd), .A(_13514_), .B(_16340_), .C(_13795_), .Y(_13796_) );
OAI21X1 OAI21X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_13792_), .B(_13793_), .C(_13483_), .Y(_13797_) );
NAND3X1 NAND3X1_3093 ( .gnd(gnd), .vdd(vdd), .A(_13482_), .B(_13786_), .C(_13790_), .Y(_13798_) );
NAND3X1 NAND3X1_3094 ( .gnd(gnd), .vdd(vdd), .A(_16340_), .B(_13798_), .C(_13797_), .Y(_13799_) );
NAND2X1 NAND2X1_1828 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_213_), .B(_13799_), .Y(_13800_) );
NAND3X1 NAND3X1_3095 ( .gnd(gnd), .vdd(vdd), .A(_13513_), .B(_13796_), .C(_13800_), .Y(_13801_) );
NOR2X1 NOR2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_213_), .B(_13799_), .Y(_13802_) );
AOI21X1 AOI21X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_16340_), .B(_13795_), .C(_13514_), .Y(_13803_) );
OAI21X1 OAI21X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_13802_), .B(_13803_), .C(_13314_), .Y(_13804_) );
NAND3X1 NAND3X1_3096 ( .gnd(gnd), .vdd(vdd), .A(_13801_), .B(_13512_), .C(_13804_), .Y(_13805_) );
OAI21X1 OAI21X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_13316_), .B(_16795_), .C(_13320_), .Y(_13806_) );
OAI21X1 OAI21X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_13802_), .B(_13803_), .C(_13513_), .Y(_13807_) );
NAND3X1 NAND3X1_3097 ( .gnd(gnd), .vdd(vdd), .A(_13314_), .B(_13796_), .C(_13800_), .Y(_13808_) );
NAND3X1 NAND3X1_3098 ( .gnd(gnd), .vdd(vdd), .A(_13808_), .B(_13806_), .C(_13807_), .Y(_13809_) );
NAND3X1 NAND3X1_3099 ( .gnd(gnd), .vdd(vdd), .A(_13491_), .B(_13805_), .C(_13809_), .Y(_13810_) );
AOI21X1 AOI21X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_13808_), .B(_13807_), .C(_13806_), .Y(_13811_) );
AOI21X1 AOI21X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_13801_), .B(_13804_), .C(_13512_), .Y(_13812_) );
OAI21X1 OAI21X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_13811_), .B(_13812_), .C(_13490_), .Y(_13813_) );
NAND2X1 NAND2X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_13810_), .B(_13813_), .Y(_13814_) );
NAND3X1 NAND3X1_3100 ( .gnd(gnd), .vdd(vdd), .A(_13511_), .B(_16349_), .C(_13814_), .Y(_13815_) );
OAI21X1 OAI21X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_13811_), .B(_13812_), .C(_13491_), .Y(_13816_) );
NAND3X1 NAND3X1_3101 ( .gnd(gnd), .vdd(vdd), .A(_13490_), .B(_13805_), .C(_13809_), .Y(_13817_) );
NAND3X1 NAND3X1_3102 ( .gnd(gnd), .vdd(vdd), .A(_16349_), .B(_13817_), .C(_13816_), .Y(_13818_) );
NAND2X1 NAND2X1_1830 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_229_), .B(_13818_), .Y(_13819_) );
NAND3X1 NAND3X1_3103 ( .gnd(gnd), .vdd(vdd), .A(_13510_), .B(_13815_), .C(_13819_), .Y(_13820_) );
NOR2X1 NOR2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_229_), .B(_13818_), .Y(_13821_) );
AOI21X1 AOI21X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_16349_), .B(_13814_), .C(_13511_), .Y(_13822_) );
OAI21X1 OAI21X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_13821_), .B(_13822_), .C(_13341_), .Y(_13823_) );
NAND3X1 NAND3X1_3104 ( .gnd(gnd), .vdd(vdd), .A(_13509_), .B(_13820_), .C(_13823_), .Y(_13824_) );
OAI21X1 OAI21X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_16793_), .B(_13343_), .C(_13346_), .Y(_13825_) );
OAI21X1 OAI21X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_13821_), .B(_13822_), .C(_13510_), .Y(_13826_) );
NAND3X1 NAND3X1_3105 ( .gnd(gnd), .vdd(vdd), .A(_13341_), .B(_13815_), .C(_13819_), .Y(_13827_) );
NAND3X1 NAND3X1_3106 ( .gnd(gnd), .vdd(vdd), .A(_13825_), .B(_13827_), .C(_13826_), .Y(_13828_) );
NAND3X1 NAND3X1_3107 ( .gnd(gnd), .vdd(vdd), .A(_13498_), .B(_13824_), .C(_13828_), .Y(_13829_) );
NAND2X1 NAND2X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_13824_), .B(_13828_), .Y(_13830_) );
AOI21X1 AOI21X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_13499_), .B(_13830_), .C(_16546_), .Y(_13831_) );
NAND3X1 NAND3X1_3108 ( .gnd(gnd), .vdd(vdd), .A(_13508_), .B(_13829_), .C(_13831_), .Y(_13832_) );
AOI21X1 AOI21X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_13827_), .B(_13826_), .C(_13825_), .Y(_13833_) );
AOI21X1 AOI21X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_13820_), .B(_13823_), .C(_13509_), .Y(_13834_) );
OAI21X1 OAI21X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_13833_), .B(_13834_), .C(_13499_), .Y(_13835_) );
NAND3X1 NAND3X1_3109 ( .gnd(gnd), .vdd(vdd), .A(_16357_), .B(_13829_), .C(_13835_), .Y(_13836_) );
NAND2X1 NAND2X1_1832 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_245_), .B(_13836_), .Y(_13837_) );
NAND3X1 NAND3X1_3110 ( .gnd(gnd), .vdd(vdd), .A(_13358_), .B(_13832_), .C(_13837_), .Y(_13838_) );
INVX1 INVX1_1946 ( .gnd(gnd), .vdd(vdd), .A(_13358_), .Y(_13839_) );
NOR2X1 NOR2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_245_), .B(_13836_), .Y(_13840_) );
AOI21X1 AOI21X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_13829_), .B(_13831_), .C(_13508_), .Y(_13841_) );
OAI21X1 OAI21X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_13840_), .B(_13841_), .C(_13839_), .Y(_13842_) );
NAND3X1 NAND3X1_3111 ( .gnd(gnd), .vdd(vdd), .A(_13838_), .B(_13507_), .C(_13842_), .Y(_13843_) );
AOI21X1 AOI21X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_13366_), .B(_16791_), .C(_13370_), .Y(_13844_) );
NOR3X1 NOR3X1_407 ( .gnd(gnd), .vdd(vdd), .A(_13839_), .B(_13841_), .C(_13840_), .Y(_13845_) );
AOI21X1 AOI21X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_13832_), .B(_13837_), .C(_13358_), .Y(_13846_) );
OAI21X1 OAI21X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_13845_), .B(_13846_), .C(_13844_), .Y(_13847_) );
NAND3X1 NAND3X1_3112 ( .gnd(gnd), .vdd(vdd), .A(_13506_), .B(_13843_), .C(_13847_), .Y(_13848_) );
INVX1 INVX1_1947 ( .gnd(gnd), .vdd(vdd), .A(_13506_), .Y(_13849_) );
NAND3X1 NAND3X1_3113 ( .gnd(gnd), .vdd(vdd), .A(_13838_), .B(_13844_), .C(_13842_), .Y(_13850_) );
OAI21X1 OAI21X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_13845_), .B(_13846_), .C(_13507_), .Y(_13851_) );
NAND3X1 NAND3X1_3114 ( .gnd(gnd), .vdd(vdd), .A(_13849_), .B(_13850_), .C(_13851_), .Y(_13852_) );
NAND2X1 NAND2X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_13848_), .B(_13852_), .Y(_13853_) );
XNOR2X1 XNOR2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_13853_), .B(_13382_), .Y(module_3_H_5_) );
AOI21X1 AOI21X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_13848_), .B(_13852_), .C(_13382_), .Y(_13854_) );
AOI21X1 AOI21X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_13838_), .B(_13507_), .C(_13846_), .Y(_13855_) );
AOI21X1 AOI21X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_13815_), .B(_13819_), .C(_13341_), .Y(_13856_) );
AOI21X1 AOI21X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_13827_), .B(_13825_), .C(_13856_), .Y(_13857_) );
INVX1 INVX1_1948 ( .gnd(gnd), .vdd(vdd), .A(_16527_), .Y(_13858_) );
INVX1 INVX1_1949 ( .gnd(gnd), .vdd(vdd), .A(_16528_), .Y(_13859_) );
NOR2X1 NOR2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_13859_), .B(_13858_), .Y(_13860_) );
INVX1 INVX1_1950 ( .gnd(gnd), .vdd(vdd), .A(_13860_), .Y(_13861_) );
AOI21X1 AOI21X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_13796_), .B(_13800_), .C(_13314_), .Y(_13862_) );
AOI21X1 AOI21X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_13808_), .B(_13806_), .C(_13862_), .Y(_13863_) );
INVX1 INVX1_1951 ( .gnd(gnd), .vdd(vdd), .A(_16517_), .Y(_13864_) );
AOI21X1 AOI21X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_13777_), .B(_13781_), .C(_13293_), .Y(_13865_) );
AOI21X1 AOI21X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_13789_), .B(_13787_), .C(_13865_), .Y(_13866_) );
NOR2X1 NOR2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_16507_), .B(_16506_), .Y(_13867_) );
INVX2 INVX2_487 ( .gnd(gnd), .vdd(vdd), .A(_13867_), .Y(_13868_) );
NOR3X1 NOR3X1_408 ( .gnd(gnd), .vdd(vdd), .A(_13519_), .B(_13765_), .C(_13764_), .Y(_13869_) );
OAI21X1 OAI21X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_13869_), .B(_13518_), .C(_13769_), .Y(_13870_) );
INVX2 INVX2_488 ( .gnd(gnd), .vdd(vdd), .A(_16499_), .Y(_13871_) );
AOI21X1 AOI21X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_13740_), .B(_13744_), .C(_13249_), .Y(_13872_) );
AOI21X1 AOI21X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_13752_), .B(_13750_), .C(_13872_), .Y(_13873_) );
INVX1 INVX1_1952 ( .gnd(gnd), .vdd(vdd), .A(_13732_), .Y(_13874_) );
AOI21X1 AOI21X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_13733_), .B(_13731_), .C(_13874_), .Y(_13875_) );
NOR2X1 NOR2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_16478_), .B(_16479_), .Y(_13876_) );
INVX1 INVX1_1953 ( .gnd(gnd), .vdd(vdd), .A(_13876_), .Y(_13877_) );
OAI21X1 OAI21X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_13706_), .B(_13528_), .C(_13713_), .Y(_13878_) );
INVX2 INVX2_489 ( .gnd(gnd), .vdd(vdd), .A(_13704_), .Y(_13879_) );
AOI21X1 AOI21X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_13681_), .B(_13677_), .C(_13172_), .Y(_13880_) );
OAI21X1 OAI21X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_13880_), .B(_13530_), .C(_13689_), .Y(_13881_) );
INVX2 INVX2_490 ( .gnd(gnd), .vdd(vdd), .A(_13677_), .Y(_13882_) );
NAND2X1 NAND2X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_13661_), .B(_13674_), .Y(_13883_) );
INVX2 INVX2_491 ( .gnd(gnd), .vdd(vdd), .A(_13656_), .Y(_13884_) );
NAND2X1 NAND2X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_13647_), .B(_13649_), .Y(_13885_) );
INVX2 INVX2_492 ( .gnd(gnd), .vdd(vdd), .A(_13635_), .Y(_13886_) );
NAND2X1 NAND2X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_13626_), .B(_13628_), .Y(_13887_) );
INVX2 INVX2_493 ( .gnd(gnd), .vdd(vdd), .A(_13614_), .Y(_13888_) );
NAND2X1 NAND2X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_13604_), .B(_13606_), .Y(_13889_) );
INVX2 INVX2_494 ( .gnd(gnd), .vdd(vdd), .A(_13592_), .Y(_13890_) );
INVX1 INVX1_1954 ( .gnd(gnd), .vdd(vdd), .A(_13584_), .Y(_13891_) );
OAI21X1 OAI21X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_13891_), .B(_13540_), .C(_13583_), .Y(_13892_) );
INVX2 INVX2_495 ( .gnd(gnd), .vdd(vdd), .A(_13572_), .Y(_13893_) );
NAND3X1 NAND3X1_3115 ( .gnd(gnd), .vdd(vdd), .A(_16835_), .B(_13552_), .C(_13556_), .Y(_13894_) );
INVX1 INVX1_1955 ( .gnd(gnd), .vdd(vdd), .A(_13552_), .Y(_13895_) );
NAND2X1 NAND2X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_16374_), .B(_16378_), .Y(_13896_) );
INVX1 INVX1_1956 ( .gnd(gnd), .vdd(vdd), .A(_13896_), .Y(_13897_) );
INVX1 INVX1_1957 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_6_), .Y(_13898_) );
AND2X2 AND2X2_311 ( .gnd(gnd), .vdd(vdd), .A(_13549_), .B(_13898_), .Y(_13899_) );
NOR2X1 NOR2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_13898_), .B(_13549_), .Y(_13900_) );
OAI21X1 OAI21X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_13899_), .B(_13900_), .C(_13897_), .Y(_13901_) );
NOR2X1 NOR2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_13900_), .B(_13899_), .Y(_13902_) );
OAI21X1 OAI21X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_16375_), .B(_16376_), .C(_13902_), .Y(_13903_) );
NAND3X1 NAND3X1_3116 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_22_), .B(_13901_), .C(_13903_), .Y(_13904_) );
INVX1 INVX1_1958 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_22_), .Y(_13905_) );
OAI21X1 OAI21X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_13899_), .B(_13900_), .C(_13896_), .Y(_13906_) );
NAND2X1 NAND2X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_13897_), .B(_13902_), .Y(_13907_) );
NAND3X1 NAND3X1_3117 ( .gnd(gnd), .vdd(vdd), .A(_13905_), .B(_13906_), .C(_13907_), .Y(_13908_) );
NAND3X1 NAND3X1_3118 ( .gnd(gnd), .vdd(vdd), .A(_13895_), .B(_13908_), .C(_13904_), .Y(_13909_) );
AOI21X1 AOI21X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_13906_), .B(_13907_), .C(_13905_), .Y(_13910_) );
AOI21X1 AOI21X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_13901_), .B(_13903_), .C(module_3_W_22_), .Y(_13911_) );
OAI21X1 OAI21X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_13911_), .B(_13910_), .C(_13552_), .Y(_13912_) );
NAND2X1 NAND2X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_13909_), .B(_13912_), .Y(_13913_) );
AOI21X1 AOI21X1_1958 ( .gnd(gnd), .vdd(vdd), .A(_13894_), .B(_13564_), .C(_13913_), .Y(_13914_) );
INVX1 INVX1_1959 ( .gnd(gnd), .vdd(vdd), .A(_13914_), .Y(_13915_) );
OAI21X1 OAI21X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_13542_), .B(_13561_), .C(_13894_), .Y(_13916_) );
INVX1 INVX1_1960 ( .gnd(gnd), .vdd(vdd), .A(_13913_), .Y(_13917_) );
OR2X2 OR2X2_342 ( .gnd(gnd), .vdd(vdd), .A(_13917_), .B(_13916_), .Y(_13918_) );
INVX2 INVX2_496 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_10_), .Y(_13919_) );
NOR2X1 NOR2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_16387_), .B(_16385_), .Y(_13920_) );
XNOR2X1 XNOR2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_13920_), .B(_13919_), .Y(_13921_) );
NAND3X1 NAND3X1_3119 ( .gnd(gnd), .vdd(vdd), .A(_13915_), .B(_13921_), .C(_13918_), .Y(_13922_) );
NOR2X1 NOR2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_13916_), .B(_13917_), .Y(_13923_) );
INVX1 INVX1_1961 ( .gnd(gnd), .vdd(vdd), .A(_13921_), .Y(_13924_) );
OAI21X1 OAI21X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_13923_), .B(_13914_), .C(_13924_), .Y(_13925_) );
NAND3X1 NAND3X1_3120 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf3_), .B(_13925_), .C(_13922_), .Y(_13926_) );
INVX2 INVX2_497 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf2_), .Y(_13927_) );
NAND3X1 NAND3X1_3121 ( .gnd(gnd), .vdd(vdd), .A(_13915_), .B(_13924_), .C(_13918_), .Y(_13928_) );
OAI21X1 OAI21X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_13923_), .B(_13914_), .C(_13921_), .Y(_13929_) );
NAND3X1 NAND3X1_3122 ( .gnd(gnd), .vdd(vdd), .A(_13927_), .B(_13929_), .C(_13928_), .Y(_13930_) );
NAND3X1 NAND3X1_3123 ( .gnd(gnd), .vdd(vdd), .A(_13893_), .B(_13926_), .C(_13930_), .Y(_13931_) );
NAND3X1 NAND3X1_3124 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf1_), .B(_13929_), .C(_13928_), .Y(_13932_) );
NAND3X1 NAND3X1_3125 ( .gnd(gnd), .vdd(vdd), .A(_13927_), .B(_13925_), .C(_13922_), .Y(_13933_) );
NAND3X1 NAND3X1_3126 ( .gnd(gnd), .vdd(vdd), .A(_13572_), .B(_13932_), .C(_13933_), .Y(_13934_) );
NAND3X1 NAND3X1_3127 ( .gnd(gnd), .vdd(vdd), .A(_13892_), .B(_13931_), .C(_13934_), .Y(_13935_) );
INVX1 INVX1_1962 ( .gnd(gnd), .vdd(vdd), .A(_13583_), .Y(_13936_) );
NOR2X1 NOR2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_13936_), .B(_13590_), .Y(_13937_) );
AOI21X1 AOI21X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_13932_), .B(_13933_), .C(_13572_), .Y(_13938_) );
AOI21X1 AOI21X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_13926_), .B(_13930_), .C(_13893_), .Y(_13939_) );
OAI21X1 OAI21X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_13938_), .B(_13939_), .C(_13937_), .Y(_13940_) );
NOR2X1 NOR2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_16397_), .B(_16404_), .Y(_13941_) );
NAND2X1 NAND2X1_1841 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_26_), .B(module_3_W_10_), .Y(_13942_) );
INVX1 INVX1_1963 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_26_), .Y(_13943_) );
NAND2X1 NAND2X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_13943_), .B(_13919_), .Y(_13944_) );
AND2X2 AND2X2_312 ( .gnd(gnd), .vdd(vdd), .A(_13944_), .B(_13942_), .Y(_13945_) );
NAND2X1 NAND2X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_13402_), .B(_13945_), .Y(_13946_) );
NAND2X1 NAND2X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_13942_), .B(_13944_), .Y(_13947_) );
OAI21X1 OAI21X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_13400_), .B(_13401_), .C(_13947_), .Y(_13948_) );
NAND3X1 NAND3X1_3128 ( .gnd(gnd), .vdd(vdd), .A(_13946_), .B(_13948_), .C(_13406_), .Y(_13949_) );
OAI21X1 OAI21X1_2192 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_24_), .B(module_3_W_8_), .C(_13404_), .Y(_13950_) );
INVX1 INVX1_1964 ( .gnd(gnd), .vdd(vdd), .A(_13402_), .Y(_13951_) );
NOR2X1 NOR2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_13951_), .B(_13947_), .Y(_13952_) );
NOR2X1 NOR2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_13402_), .B(_13945_), .Y(_13953_) );
OAI21X1 OAI21X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_13953_), .B(_13952_), .C(_13950_), .Y(_13954_) );
NAND2X1 NAND2X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_13954_), .B(_13949_), .Y(_13955_) );
XNOR2X1 XNOR2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_13941_), .B(_13955_), .Y(_13956_) );
NAND3X1 NAND3X1_3129 ( .gnd(gnd), .vdd(vdd), .A(_13935_), .B(_13956_), .C(_13940_), .Y(_13957_) );
NAND3X1 NAND3X1_3130 ( .gnd(gnd), .vdd(vdd), .A(_13572_), .B(_13926_), .C(_13930_), .Y(_13958_) );
NAND3X1 NAND3X1_3131 ( .gnd(gnd), .vdd(vdd), .A(_13893_), .B(_13932_), .C(_13933_), .Y(_13959_) );
AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_13583_), .B(_13585_), .C(_13958_), .D(_13959_), .Y(_13960_) );
AOI21X1 AOI21X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_13931_), .B(_13934_), .C(_13892_), .Y(_13961_) );
INVX1 INVX1_1965 ( .gnd(gnd), .vdd(vdd), .A(_13956_), .Y(_13962_) );
OAI21X1 OAI21X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_13960_), .B(_13961_), .C(_13962_), .Y(_13963_) );
NAND3X1 NAND3X1_3132 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf3_), .B(_13957_), .C(_13963_), .Y(_13964_) );
INVX1 INVX1_1966 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf2_), .Y(_13965_) );
NAND3X1 NAND3X1_3133 ( .gnd(gnd), .vdd(vdd), .A(_13935_), .B(_13962_), .C(_13940_), .Y(_13966_) );
OAI21X1 OAI21X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_13960_), .B(_13961_), .C(_13956_), .Y(_13967_) );
NAND3X1 NAND3X1_3134 ( .gnd(gnd), .vdd(vdd), .A(_13965_), .B(_13966_), .C(_13967_), .Y(_13968_) );
NAND3X1 NAND3X1_3135 ( .gnd(gnd), .vdd(vdd), .A(_13890_), .B(_13964_), .C(_13968_), .Y(_13969_) );
NAND3X1 NAND3X1_3136 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf1_), .B(_13966_), .C(_13967_), .Y(_13970_) );
NAND3X1 NAND3X1_3137 ( .gnd(gnd), .vdd(vdd), .A(_13965_), .B(_13957_), .C(_13963_), .Y(_13971_) );
NAND3X1 NAND3X1_3138 ( .gnd(gnd), .vdd(vdd), .A(_13592_), .B(_13970_), .C(_13971_), .Y(_13972_) );
NAND3X1 NAND3X1_3139 ( .gnd(gnd), .vdd(vdd), .A(_13969_), .B(_13972_), .C(_13889_), .Y(_13973_) );
AND2X2 AND2X2_313 ( .gnd(gnd), .vdd(vdd), .A(_13606_), .B(_13604_), .Y(_13974_) );
AOI21X1 AOI21X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_13970_), .B(_13971_), .C(_13592_), .Y(_13975_) );
AOI21X1 AOI21X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_13964_), .B(_13968_), .C(_13890_), .Y(_13976_) );
OAI21X1 OAI21X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_13975_), .B(_13976_), .C(_13974_), .Y(_13977_) );
NOR2X1 NOR2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_16414_), .B(_16411_), .Y(_13978_) );
NOR2X1 NOR2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_13399_), .B(_13413_), .Y(_13979_) );
INVX1 INVX1_1967 ( .gnd(gnd), .vdd(vdd), .A(_13411_), .Y(_13980_) );
INVX1 INVX1_1968 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .Y(_13981_) );
NAND2X1 NAND2X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_13981_), .B(_13955_), .Y(_13982_) );
NAND3X1 NAND3X1_3140 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .B(_13954_), .C(_13949_), .Y(_13983_) );
NAND2X1 NAND2X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_13983_), .B(_13982_), .Y(_13984_) );
NOR2X1 NOR2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_13980_), .B(_13984_), .Y(_13985_) );
AOI21X1 AOI21X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_13983_), .B(_13982_), .C(_13411_), .Y(_13986_) );
NOR2X1 NOR2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_13986_), .B(_13985_), .Y(_13987_) );
NAND2X1 NAND2X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_13979_), .B(_13987_), .Y(_13988_) );
OAI21X1 OAI21X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_13985_), .B(_13986_), .C(_13414_), .Y(_13989_) );
NAND2X1 NAND2X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_13989_), .B(_13988_), .Y(_13990_) );
XNOR2X1 XNOR2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_13978_), .B(_13990_), .Y(_13991_) );
NAND3X1 NAND3X1_3141 ( .gnd(gnd), .vdd(vdd), .A(_13973_), .B(_13991_), .C(_13977_), .Y(_13992_) );
NAND3X1 NAND3X1_3142 ( .gnd(gnd), .vdd(vdd), .A(_13592_), .B(_13964_), .C(_13968_), .Y(_13993_) );
NAND3X1 NAND3X1_3143 ( .gnd(gnd), .vdd(vdd), .A(_13890_), .B(_13970_), .C(_13971_), .Y(_13994_) );
AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_13604_), .B(_13606_), .C(_13993_), .D(_13994_), .Y(_13995_) );
AOI21X1 AOI21X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_13969_), .B(_13972_), .C(_13889_), .Y(_13996_) );
INVX1 INVX1_1969 ( .gnd(gnd), .vdd(vdd), .A(_13991_), .Y(_13997_) );
OAI21X1 OAI21X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_13995_), .B(_13996_), .C(_13997_), .Y(_13998_) );
NAND3X1 NAND3X1_3144 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf0_), .B(_13998_), .C(_13992_), .Y(_13999_) );
INVX1 INVX1_1970 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf3_), .Y(_14000_) );
NAND3X1 NAND3X1_3145 ( .gnd(gnd), .vdd(vdd), .A(_13973_), .B(_13997_), .C(_13977_), .Y(_14001_) );
OAI21X1 OAI21X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_13995_), .B(_13996_), .C(_13991_), .Y(_14002_) );
NAND3X1 NAND3X1_3146 ( .gnd(gnd), .vdd(vdd), .A(_14000_), .B(_14002_), .C(_14001_), .Y(_14003_) );
NAND3X1 NAND3X1_3147 ( .gnd(gnd), .vdd(vdd), .A(_13888_), .B(_13999_), .C(_14003_), .Y(_14004_) );
NAND3X1 NAND3X1_3148 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf2_), .B(_14002_), .C(_14001_), .Y(_14005_) );
NAND3X1 NAND3X1_3149 ( .gnd(gnd), .vdd(vdd), .A(_14000_), .B(_13998_), .C(_13992_), .Y(_14006_) );
NAND3X1 NAND3X1_3150 ( .gnd(gnd), .vdd(vdd), .A(_13614_), .B(_14005_), .C(_14006_), .Y(_14007_) );
NAND3X1 NAND3X1_3151 ( .gnd(gnd), .vdd(vdd), .A(_14004_), .B(_14007_), .C(_13887_), .Y(_14008_) );
AND2X2 AND2X2_314 ( .gnd(gnd), .vdd(vdd), .A(_13628_), .B(_13626_), .Y(_14009_) );
AOI21X1 AOI21X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_14005_), .B(_14006_), .C(_13614_), .Y(_14010_) );
AOI21X1 AOI21X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_13999_), .B(_14003_), .C(_13888_), .Y(_14011_) );
OAI21X1 OAI21X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_14010_), .B(_14011_), .C(_14009_), .Y(_14012_) );
INVX2 INVX2_498 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf3_), .Y(_14013_) );
AND2X2 AND2X2_315 ( .gnd(gnd), .vdd(vdd), .A(_13987_), .B(_13979_), .Y(_14014_) );
INVX1 INVX1_1971 ( .gnd(gnd), .vdd(vdd), .A(_13989_), .Y(_14015_) );
OAI21X1 OAI21X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_14014_), .B(_14015_), .C(_14013_), .Y(_14016_) );
OR2X2 OR2X2_343 ( .gnd(gnd), .vdd(vdd), .A(_13990_), .B(_14013_), .Y(_14017_) );
NAND3X1 NAND3X1_3152 ( .gnd(gnd), .vdd(vdd), .A(_13417_), .B(_14016_), .C(_14017_), .Y(_14018_) );
INVX1 INVX1_1972 ( .gnd(gnd), .vdd(vdd), .A(_13417_), .Y(_14019_) );
INVX1 INVX1_1973 ( .gnd(gnd), .vdd(vdd), .A(_14016_), .Y(_14020_) );
NOR2X1 NOR2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_14013_), .B(_13990_), .Y(_14021_) );
OAI21X1 OAI21X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_14020_), .B(_14021_), .C(_14019_), .Y(_14022_) );
NAND2X1 NAND2X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_14018_), .B(_14022_), .Y(_14023_) );
OR2X2 OR2X2_344 ( .gnd(gnd), .vdd(vdd), .A(_14023_), .B(_13420_), .Y(_14024_) );
NOR3X1 NOR3X1_409 ( .gnd(gnd), .vdd(vdd), .A(_14019_), .B(_14021_), .C(_14020_), .Y(_14025_) );
AOI21X1 AOI21X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_14016_), .B(_14017_), .C(_13417_), .Y(_14026_) );
OAI21X1 OAI21X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_14025_), .B(_14026_), .C(_13420_), .Y(_14027_) );
NAND2X1 NAND2X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_14027_), .B(_14024_), .Y(_14028_) );
XNOR2X1 XNOR2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_16643_), .B(_14028_), .Y(_14029_) );
NAND3X1 NAND3X1_3153 ( .gnd(gnd), .vdd(vdd), .A(_14008_), .B(_14029_), .C(_14012_), .Y(_14030_) );
NAND3X1 NAND3X1_3154 ( .gnd(gnd), .vdd(vdd), .A(_13614_), .B(_13999_), .C(_14003_), .Y(_14031_) );
NAND3X1 NAND3X1_3155 ( .gnd(gnd), .vdd(vdd), .A(_13888_), .B(_14005_), .C(_14006_), .Y(_14032_) );
AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_13626_), .B(_13628_), .C(_14031_), .D(_14032_), .Y(_14033_) );
AOI21X1 AOI21X1_1969 ( .gnd(gnd), .vdd(vdd), .A(_14004_), .B(_14007_), .C(_13887_), .Y(_14034_) );
INVX1 INVX1_1974 ( .gnd(gnd), .vdd(vdd), .A(_14029_), .Y(_14035_) );
OAI21X1 OAI21X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_14033_), .B(_14034_), .C(_14035_), .Y(_14036_) );
NAND3X1 NAND3X1_3156 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf0_), .B(_14030_), .C(_14036_), .Y(_14037_) );
INVX1 INVX1_1975 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf3_), .Y(_14038_) );
OAI21X1 OAI21X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_14033_), .B(_14034_), .C(_14029_), .Y(_14039_) );
NAND3X1 NAND3X1_3157 ( .gnd(gnd), .vdd(vdd), .A(_14008_), .B(_14035_), .C(_14012_), .Y(_14040_) );
NAND3X1 NAND3X1_3158 ( .gnd(gnd), .vdd(vdd), .A(_14038_), .B(_14040_), .C(_14039_), .Y(_14041_) );
NAND3X1 NAND3X1_3159 ( .gnd(gnd), .vdd(vdd), .A(_13886_), .B(_14037_), .C(_14041_), .Y(_14042_) );
NAND3X1 NAND3X1_3160 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf2_), .B(_14040_), .C(_14039_), .Y(_14043_) );
NAND3X1 NAND3X1_3161 ( .gnd(gnd), .vdd(vdd), .A(_14038_), .B(_14030_), .C(_14036_), .Y(_14044_) );
NAND3X1 NAND3X1_3162 ( .gnd(gnd), .vdd(vdd), .A(_13635_), .B(_14043_), .C(_14044_), .Y(_14045_) );
NAND3X1 NAND3X1_3163 ( .gnd(gnd), .vdd(vdd), .A(_14042_), .B(_14045_), .C(_13885_), .Y(_14046_) );
AND2X2 AND2X2_316 ( .gnd(gnd), .vdd(vdd), .A(_13649_), .B(_13647_), .Y(_14047_) );
AOI21X1 AOI21X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_14043_), .B(_14044_), .C(_13635_), .Y(_14048_) );
AOI21X1 AOI21X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_14037_), .B(_14041_), .C(_13886_), .Y(_14049_) );
OAI21X1 OAI21X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_14048_), .B(_14049_), .C(_14047_), .Y(_14050_) );
INVX1 INVX1_1976 ( .gnd(gnd), .vdd(vdd), .A(_13425_), .Y(_14051_) );
INVX1 INVX1_1977 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf0_), .Y(_14052_) );
NOR2X1 NOR2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_13420_), .B(_14023_), .Y(_14053_) );
INVX1 INVX1_1978 ( .gnd(gnd), .vdd(vdd), .A(_14027_), .Y(_14054_) );
OAI21X1 OAI21X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_14054_), .B(_14053_), .C(_14052_), .Y(_14055_) );
INVX1 INVX1_1979 ( .gnd(gnd), .vdd(vdd), .A(_14055_), .Y(_14056_) );
NOR2X1 NOR2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_14052_), .B(_14028_), .Y(_14057_) );
NOR3X1 NOR3X1_410 ( .gnd(gnd), .vdd(vdd), .A(_14056_), .B(_14051_), .C(_14057_), .Y(_14058_) );
NOR2X1 NOR2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_14053_), .B(_14054_), .Y(_14059_) );
NAND2X1 NAND2X1_1852 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf3_), .B(_14059_), .Y(_14060_) );
AOI21X1 AOI21X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_14055_), .B(_14060_), .C(_13425_), .Y(_14061_) );
NOR3X1 NOR3X1_411 ( .gnd(gnd), .vdd(vdd), .A(_13428_), .B(_14061_), .C(_14058_), .Y(_14062_) );
INVX2 INVX2_499 ( .gnd(gnd), .vdd(vdd), .A(_13428_), .Y(_14063_) );
NAND3X1 NAND3X1_3164 ( .gnd(gnd), .vdd(vdd), .A(_13425_), .B(_14055_), .C(_14060_), .Y(_14064_) );
OAI21X1 OAI21X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_14057_), .B(_14056_), .C(_14051_), .Y(_14065_) );
AOI21X1 AOI21X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_14064_), .B(_14065_), .C(_14063_), .Y(_14066_) );
NOR2X1 NOR2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_14066_), .B(_14062_), .Y(_14067_) );
OAI21X1 OAI21X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_16434_), .B(_16435_), .C(_14067_), .Y(_14068_) );
NOR2X1 NOR2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_16435_), .B(_16434_), .Y(_14069_) );
OAI21X1 OAI21X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_14062_), .B(_14066_), .C(_14069_), .Y(_14070_) );
NAND2X1 NAND2X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_14068_), .B(_14070_), .Y(_14071_) );
NAND3X1 NAND3X1_3165 ( .gnd(gnd), .vdd(vdd), .A(_14046_), .B(_14071_), .C(_14050_), .Y(_14072_) );
NAND3X1 NAND3X1_3166 ( .gnd(gnd), .vdd(vdd), .A(_13635_), .B(_14037_), .C(_14041_), .Y(_14073_) );
NAND3X1 NAND3X1_3167 ( .gnd(gnd), .vdd(vdd), .A(_13886_), .B(_14043_), .C(_14044_), .Y(_14074_) );
AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_13647_), .B(_13649_), .C(_14073_), .D(_14074_), .Y(_14075_) );
AOI21X1 AOI21X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_14042_), .B(_14045_), .C(_13885_), .Y(_14076_) );
INVX1 INVX1_1980 ( .gnd(gnd), .vdd(vdd), .A(_14071_), .Y(_14077_) );
OAI21X1 OAI21X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_14075_), .B(_14076_), .C(_14077_), .Y(_14078_) );
NAND3X1 NAND3X1_3168 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf0_), .B(_14072_), .C(_14078_), .Y(_14079_) );
INVX1 INVX1_1981 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf3_), .Y(_14080_) );
OAI21X1 OAI21X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_14075_), .B(_14076_), .C(_14071_), .Y(_14081_) );
NAND3X1 NAND3X1_3169 ( .gnd(gnd), .vdd(vdd), .A(_14046_), .B(_14077_), .C(_14050_), .Y(_14082_) );
NAND3X1 NAND3X1_3170 ( .gnd(gnd), .vdd(vdd), .A(_14080_), .B(_14082_), .C(_14081_), .Y(_14083_) );
NAND3X1 NAND3X1_3171 ( .gnd(gnd), .vdd(vdd), .A(_13884_), .B(_14079_), .C(_14083_), .Y(_14084_) );
NAND3X1 NAND3X1_3172 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf2_), .B(_14082_), .C(_14081_), .Y(_14085_) );
NAND3X1 NAND3X1_3173 ( .gnd(gnd), .vdd(vdd), .A(_14080_), .B(_14072_), .C(_14078_), .Y(_14086_) );
NAND3X1 NAND3X1_3174 ( .gnd(gnd), .vdd(vdd), .A(_13656_), .B(_14085_), .C(_14086_), .Y(_14087_) );
NAND3X1 NAND3X1_3175 ( .gnd(gnd), .vdd(vdd), .A(_14084_), .B(_14087_), .C(_13883_), .Y(_14088_) );
AND2X2 AND2X2_317 ( .gnd(gnd), .vdd(vdd), .A(_13674_), .B(_13661_), .Y(_14089_) );
AOI21X1 AOI21X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_14085_), .B(_14086_), .C(_13656_), .Y(_14090_) );
AOI21X1 AOI21X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_14079_), .B(_14083_), .C(_13884_), .Y(_14091_) );
OAI21X1 OAI21X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_14090_), .B(_14091_), .C(_14089_), .Y(_14092_) );
INVX1 INVX1_1982 ( .gnd(gnd), .vdd(vdd), .A(_13433_), .Y(_14093_) );
NAND3X1 NAND3X1_3176 ( .gnd(gnd), .vdd(vdd), .A(_14064_), .B(_14065_), .C(_14063_), .Y(_14094_) );
OAI21X1 OAI21X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_14058_), .B(_14061_), .C(_13428_), .Y(_14095_) );
AOI21X1 AOI21X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_14094_), .B(_14095_), .C(bloque_datos_58_bF_buf1_), .Y(_14096_) );
INVX1 INVX1_1983 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf0_), .Y(_14097_) );
NOR3X1 NOR3X1_412 ( .gnd(gnd), .vdd(vdd), .A(_14097_), .B(_14066_), .C(_14062_), .Y(_14098_) );
NOR3X1 NOR3X1_413 ( .gnd(gnd), .vdd(vdd), .A(_14093_), .B(_14096_), .C(_14098_), .Y(_14099_) );
OAI21X1 OAI21X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_14062_), .B(_14066_), .C(_14097_), .Y(_14100_) );
NAND3X1 NAND3X1_3177 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf4_), .B(_14094_), .C(_14095_), .Y(_14101_) );
AOI21X1 AOI21X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_14101_), .B(_14100_), .C(_13433_), .Y(_14102_) );
NOR3X1 NOR3X1_414 ( .gnd(gnd), .vdd(vdd), .A(_13436_), .B(_14102_), .C(_14099_), .Y(_14103_) );
NOR2X1 NOR2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_13396_), .B(_13435_), .Y(_14104_) );
NAND3X1 NAND3X1_3178 ( .gnd(gnd), .vdd(vdd), .A(_13433_), .B(_14101_), .C(_14100_), .Y(_14105_) );
OAI21X1 OAI21X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_14098_), .B(_14096_), .C(_14093_), .Y(_14106_) );
AOI21X1 AOI21X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_14105_), .B(_14106_), .C(_14104_), .Y(_14107_) );
NOR2X1 NOR2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_14107_), .B(_14103_), .Y(_14108_) );
OAI21X1 OAI21X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_16454_), .B(_16455_), .C(_14108_), .Y(_14109_) );
NOR2X1 NOR2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_16455_), .B(_16454_), .Y(_14110_) );
OAI21X1 OAI21X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_14103_), .B(_14107_), .C(_14110_), .Y(_14111_) );
NAND2X1 NAND2X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_14109_), .B(_14111_), .Y(_14112_) );
NAND3X1 NAND3X1_3179 ( .gnd(gnd), .vdd(vdd), .A(_14088_), .B(_14112_), .C(_14092_), .Y(_14113_) );
NAND3X1 NAND3X1_3180 ( .gnd(gnd), .vdd(vdd), .A(_13656_), .B(_14079_), .C(_14083_), .Y(_14114_) );
NAND3X1 NAND3X1_3181 ( .gnd(gnd), .vdd(vdd), .A(_13884_), .B(_14085_), .C(_14086_), .Y(_14115_) );
AOI22X1 AOI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_13661_), .B(_13674_), .C(_14114_), .D(_14115_), .Y(_14116_) );
AOI21X1 AOI21X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_14084_), .B(_14087_), .C(_13883_), .Y(_14117_) );
INVX1 INVX1_1984 ( .gnd(gnd), .vdd(vdd), .A(_14112_), .Y(_14118_) );
OAI21X1 OAI21X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_14117_), .B(_14116_), .C(_14118_), .Y(_14119_) );
NAND3X1 NAND3X1_3182 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf1_), .B(_14119_), .C(_14113_), .Y(_14120_) );
INVX1 INVX1_1985 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf0_), .Y(_14121_) );
OAI21X1 OAI21X1_2220 ( .gnd(gnd), .vdd(vdd), .A(_14117_), .B(_14116_), .C(_14112_), .Y(_14122_) );
NAND3X1 NAND3X1_3183 ( .gnd(gnd), .vdd(vdd), .A(_14088_), .B(_14118_), .C(_14092_), .Y(_14123_) );
NAND3X1 NAND3X1_3184 ( .gnd(gnd), .vdd(vdd), .A(_14121_), .B(_14122_), .C(_14123_), .Y(_14124_) );
NAND3X1 NAND3X1_3185 ( .gnd(gnd), .vdd(vdd), .A(_13882_), .B(_14120_), .C(_14124_), .Y(_14125_) );
NAND3X1 NAND3X1_3186 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf4_), .B(_14122_), .C(_14123_), .Y(_14126_) );
NAND3X1 NAND3X1_3187 ( .gnd(gnd), .vdd(vdd), .A(_14121_), .B(_14119_), .C(_14113_), .Y(_14127_) );
NAND3X1 NAND3X1_3188 ( .gnd(gnd), .vdd(vdd), .A(_13677_), .B(_14126_), .C(_14127_), .Y(_14128_) );
NAND3X1 NAND3X1_3189 ( .gnd(gnd), .vdd(vdd), .A(_13881_), .B(_14125_), .C(_14128_), .Y(_14129_) );
INVX1 INVX1_1986 ( .gnd(gnd), .vdd(vdd), .A(_13881_), .Y(_14130_) );
AOI21X1 AOI21X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_14126_), .B(_14127_), .C(_13677_), .Y(_14131_) );
AOI21X1 AOI21X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_14120_), .B(_14124_), .C(_13882_), .Y(_14132_) );
OAI21X1 OAI21X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_14131_), .B(_14132_), .C(_14130_), .Y(_14133_) );
INVX1 INVX1_1987 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf1_), .Y(_14134_) );
OAI21X1 OAI21X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_14103_), .B(_14107_), .C(_14134_), .Y(_14135_) );
NAND3X1 NAND3X1_3190 ( .gnd(gnd), .vdd(vdd), .A(_14104_), .B(_14105_), .C(_14106_), .Y(_14136_) );
OAI21X1 OAI21X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_14099_), .B(_14102_), .C(_13436_), .Y(_14137_) );
NAND3X1 NAND3X1_3191 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf0_), .B(_14136_), .C(_14137_), .Y(_14138_) );
NAND2X1 NAND2X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_14138_), .B(_14135_), .Y(_14139_) );
NOR2X1 NOR2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_13439_), .B(_14139_), .Y(_14140_) );
INVX1 INVX1_1988 ( .gnd(gnd), .vdd(vdd), .A(_13439_), .Y(_14141_) );
AOI21X1 AOI21X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_14138_), .B(_14135_), .C(_14141_), .Y(_14142_) );
NOR3X1 NOR3X1_415 ( .gnd(gnd), .vdd(vdd), .A(_13442_), .B(_14142_), .C(_14140_), .Y(_14143_) );
NOR2X1 NOR2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_13180_), .B(_13440_), .Y(_14144_) );
NAND3X1 NAND3X1_3192 ( .gnd(gnd), .vdd(vdd), .A(_14135_), .B(_14138_), .C(_14141_), .Y(_14145_) );
INVX1 INVX1_1989 ( .gnd(gnd), .vdd(vdd), .A(_14142_), .Y(_14146_) );
AOI21X1 AOI21X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_14145_), .B(_14146_), .C(_14144_), .Y(_14147_) );
NOR2X1 NOR2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_14147_), .B(_14143_), .Y(_14148_) );
OAI21X1 OAI21X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_16466_), .B(_16467_), .C(_14148_), .Y(_14149_) );
NOR2X1 NOR2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_16467_), .B(_16466_), .Y(_14150_) );
OAI21X1 OAI21X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_14143_), .B(_14147_), .C(_14150_), .Y(_14151_) );
NAND2X1 NAND2X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_14149_), .B(_14151_), .Y(_14152_) );
NAND3X1 NAND3X1_3193 ( .gnd(gnd), .vdd(vdd), .A(_14129_), .B(_14152_), .C(_14133_), .Y(_14153_) );
NAND3X1 NAND3X1_3194 ( .gnd(gnd), .vdd(vdd), .A(_13677_), .B(_14120_), .C(_14124_), .Y(_14154_) );
NAND3X1 NAND3X1_3195 ( .gnd(gnd), .vdd(vdd), .A(_13882_), .B(_14126_), .C(_14127_), .Y(_14155_) );
AOI21X1 AOI21X1_1985 ( .gnd(gnd), .vdd(vdd), .A(_14154_), .B(_14155_), .C(_14130_), .Y(_14156_) );
AOI21X1 AOI21X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_14125_), .B(_14128_), .C(_13881_), .Y(_14157_) );
INVX1 INVX1_1990 ( .gnd(gnd), .vdd(vdd), .A(_14152_), .Y(_14158_) );
OAI21X1 OAI21X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_14156_), .B(_14157_), .C(_14158_), .Y(_14159_) );
NAND3X1 NAND3X1_3196 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_134_), .B(_14153_), .C(_14159_), .Y(_14160_) );
INVX1 INVX1_1991 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_134_), .Y(_14161_) );
NAND3X1 NAND3X1_3197 ( .gnd(gnd), .vdd(vdd), .A(_14129_), .B(_14158_), .C(_14133_), .Y(_14162_) );
OAI21X1 OAI21X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_14156_), .B(_14157_), .C(_14152_), .Y(_14163_) );
NAND3X1 NAND3X1_3198 ( .gnd(gnd), .vdd(vdd), .A(_14161_), .B(_14162_), .C(_14163_), .Y(_14164_) );
NAND3X1 NAND3X1_3199 ( .gnd(gnd), .vdd(vdd), .A(_13879_), .B(_14160_), .C(_14164_), .Y(_14165_) );
NAND3X1 NAND3X1_3200 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_134_), .B(_14162_), .C(_14163_), .Y(_14166_) );
NAND3X1 NAND3X1_3201 ( .gnd(gnd), .vdd(vdd), .A(_14161_), .B(_14153_), .C(_14159_), .Y(_14167_) );
NAND3X1 NAND3X1_3202 ( .gnd(gnd), .vdd(vdd), .A(_13704_), .B(_14166_), .C(_14167_), .Y(_14168_) );
NAND3X1 NAND3X1_3203 ( .gnd(gnd), .vdd(vdd), .A(_13878_), .B(_14165_), .C(_14168_), .Y(_14169_) );
INVX2 INVX2_500 ( .gnd(gnd), .vdd(vdd), .A(_13878_), .Y(_14170_) );
AOI21X1 AOI21X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_14166_), .B(_14167_), .C(_13704_), .Y(_14171_) );
AOI21X1 AOI21X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_14160_), .B(_14164_), .C(_13879_), .Y(_14172_) );
OAI21X1 OAI21X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_14171_), .B(_14172_), .C(_14170_), .Y(_14173_) );
INVX1 INVX1_1992 ( .gnd(gnd), .vdd(vdd), .A(_13445_), .Y(_14174_) );
INVX1 INVX1_1993 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf3_), .Y(_14175_) );
OAI21X1 OAI21X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_14143_), .B(_14147_), .C(_14175_), .Y(_14176_) );
NAND3X1 NAND3X1_3204 ( .gnd(gnd), .vdd(vdd), .A(_14144_), .B(_14145_), .C(_14146_), .Y(_14177_) );
OAI21X1 OAI21X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_14140_), .B(_14142_), .C(_13442_), .Y(_14178_) );
NAND3X1 NAND3X1_3205 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf2_), .B(_14178_), .C(_14177_), .Y(_14179_) );
NAND3X1 NAND3X1_3206 ( .gnd(gnd), .vdd(vdd), .A(_14176_), .B(_14179_), .C(_14174_), .Y(_14180_) );
AOI21X1 AOI21X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_14178_), .B(_14177_), .C(bloque_datos_90_bF_buf1_), .Y(_14181_) );
NOR3X1 NOR3X1_416 ( .gnd(gnd), .vdd(vdd), .A(_14147_), .B(_14175_), .C(_14143_), .Y(_14182_) );
OAI21X1 OAI21X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_14182_), .B(_14181_), .C(_13445_), .Y(_14183_) );
AND2X2 AND2X2_318 ( .gnd(gnd), .vdd(vdd), .A(_14183_), .B(_14180_), .Y(_14184_) );
NAND2X1 NAND2X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_13448_), .B(_14184_), .Y(_14185_) );
INVX1 INVX1_1994 ( .gnd(gnd), .vdd(vdd), .A(_14185_), .Y(_14186_) );
NOR2X1 NOR2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_13448_), .B(_14184_), .Y(_14187_) );
NOR2X1 NOR2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_14187_), .B(_14186_), .Y(_14188_) );
INVX4 INVX4_13 ( .gnd(gnd), .vdd(vdd), .A(_14188_), .Y(_14189_) );
NAND3X1 NAND3X1_3207 ( .gnd(gnd), .vdd(vdd), .A(_14169_), .B(_14189_), .C(_14173_), .Y(_14190_) );
NAND3X1 NAND3X1_3208 ( .gnd(gnd), .vdd(vdd), .A(_13704_), .B(_14160_), .C(_14164_), .Y(_14191_) );
NAND3X1 NAND3X1_3209 ( .gnd(gnd), .vdd(vdd), .A(_13879_), .B(_14166_), .C(_14167_), .Y(_14192_) );
AOI21X1 AOI21X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_14191_), .B(_14192_), .C(_14170_), .Y(_14193_) );
AOI21X1 AOI21X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_14165_), .B(_14168_), .C(_13878_), .Y(_14194_) );
OAI21X1 OAI21X1_2232 ( .gnd(gnd), .vdd(vdd), .A(_14193_), .B(_14194_), .C(_14188_), .Y(_14195_) );
NAND3X1 NAND3X1_3210 ( .gnd(gnd), .vdd(vdd), .A(_13877_), .B(_14190_), .C(_14195_), .Y(_14196_) );
NAND2X1 NAND2X1_1858 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_150_), .B(_14196_), .Y(_14197_) );
INVX2 INVX2_501 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_150_), .Y(_14198_) );
OAI21X1 OAI21X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_14193_), .B(_14194_), .C(_14189_), .Y(_14199_) );
NAND3X1 NAND3X1_3211 ( .gnd(gnd), .vdd(vdd), .A(_14169_), .B(_14188_), .C(_14173_), .Y(_14200_) );
AOI21X1 AOI21X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_14200_), .B(_14199_), .C(_13876_), .Y(_14201_) );
NAND2X1 NAND2X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_14198_), .B(_14201_), .Y(_14202_) );
NAND3X1 NAND3X1_3212 ( .gnd(gnd), .vdd(vdd), .A(_13727_), .B(_14197_), .C(_14202_), .Y(_14203_) );
NAND2X1 NAND2X1_1860 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_150_), .B(_14201_), .Y(_14204_) );
NAND2X1 NAND2X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_14198_), .B(_14196_), .Y(_14205_) );
NAND3X1 NAND3X1_3213 ( .gnd(gnd), .vdd(vdd), .A(_13721_), .B(_14205_), .C(_14204_), .Y(_14206_) );
AOI21X1 AOI21X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_14203_), .B(_14206_), .C(_13875_), .Y(_14207_) );
INVX1 INVX1_1995 ( .gnd(gnd), .vdd(vdd), .A(_13733_), .Y(_14208_) );
OAI21X1 OAI21X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_14208_), .B(_13525_), .C(_13732_), .Y(_14209_) );
NAND3X1 NAND3X1_3214 ( .gnd(gnd), .vdd(vdd), .A(_13721_), .B(_14197_), .C(_14202_), .Y(_14210_) );
NAND3X1 NAND3X1_3215 ( .gnd(gnd), .vdd(vdd), .A(_13727_), .B(_14205_), .C(_14204_), .Y(_14211_) );
AOI21X1 AOI21X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_14210_), .B(_14211_), .C(_14209_), .Y(_14212_) );
INVX1 INVX1_1996 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_138_), .Y(_14213_) );
OAI21X1 OAI21X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_14186_), .B(_14187_), .C(_14213_), .Y(_14214_) );
NAND2X1 NAND2X1_1862 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_138_), .B(_14188_), .Y(_14215_) );
NAND2X1 NAND2X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_14214_), .B(_14215_), .Y(_14216_) );
NOR2X1 NOR2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_13453_), .B(_14216_), .Y(_14217_) );
INVX1 INVX1_1997 ( .gnd(gnd), .vdd(vdd), .A(_14217_), .Y(_14218_) );
OAI21X1 OAI21X1_2236 ( .gnd(gnd), .vdd(vdd), .A(_13391_), .B(_13450_), .C(_14216_), .Y(_14219_) );
NAND3X1 NAND3X1_3216 ( .gnd(gnd), .vdd(vdd), .A(_13456_), .B(_14219_), .C(_14218_), .Y(_14220_) );
INVX1 INVX1_1998 ( .gnd(gnd), .vdd(vdd), .A(_14219_), .Y(_14221_) );
OAI21X1 OAI21X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_14221_), .B(_14217_), .C(_13457_), .Y(_14222_) );
NAND2X1 NAND2X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_14222_), .B(_14220_), .Y(_14223_) );
INVX2 INVX2_502 ( .gnd(gnd), .vdd(vdd), .A(_14223_), .Y(_14224_) );
OAI21X1 OAI21X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_14207_), .B(_14212_), .C(_14224_), .Y(_14225_) );
NAND3X1 NAND3X1_3217 ( .gnd(gnd), .vdd(vdd), .A(_14210_), .B(_14211_), .C(_14209_), .Y(_14226_) );
AOI21X1 AOI21X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_14205_), .B(_14204_), .C(_13727_), .Y(_14227_) );
AOI21X1 AOI21X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_14197_), .B(_14202_), .C(_13721_), .Y(_14228_) );
OAI21X1 OAI21X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_14227_), .B(_14228_), .C(_13875_), .Y(_14229_) );
NAND3X1 NAND3X1_3218 ( .gnd(gnd), .vdd(vdd), .A(_14223_), .B(_14226_), .C(_14229_), .Y(_14230_) );
NAND3X1 NAND3X1_3219 ( .gnd(gnd), .vdd(vdd), .A(_16702_), .B(_14230_), .C(_14225_), .Y(_14231_) );
NAND2X1 NAND2X1_1865 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_166_), .B(_14231_), .Y(_14232_) );
INVX2 INVX2_503 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_166_), .Y(_14233_) );
NAND3X1 NAND3X1_3220 ( .gnd(gnd), .vdd(vdd), .A(_14224_), .B(_14226_), .C(_14229_), .Y(_14234_) );
OAI21X1 OAI21X1_2240 ( .gnd(gnd), .vdd(vdd), .A(_14207_), .B(_14212_), .C(_14223_), .Y(_14235_) );
AOI21X1 AOI21X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_14234_), .B(_14235_), .C(_16489_), .Y(_14236_) );
NAND2X1 NAND2X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_14233_), .B(_14236_), .Y(_14237_) );
NAND3X1 NAND3X1_3221 ( .gnd(gnd), .vdd(vdd), .A(_13746_), .B(_14232_), .C(_14237_), .Y(_14238_) );
NAND2X1 NAND2X1_1867 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_166_), .B(_14236_), .Y(_14239_) );
NAND2X1 NAND2X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_14233_), .B(_14231_), .Y(_14240_) );
NAND3X1 NAND3X1_3222 ( .gnd(gnd), .vdd(vdd), .A(_13740_), .B(_14240_), .C(_14239_), .Y(_14241_) );
AOI21X1 AOI21X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_14238_), .B(_14241_), .C(_13873_), .Y(_14242_) );
NOR3X1 NOR3X1_417 ( .gnd(gnd), .vdd(vdd), .A(_13747_), .B(_13522_), .C(_13746_), .Y(_14243_) );
OAI21X1 OAI21X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_14243_), .B(_13521_), .C(_13751_), .Y(_14244_) );
NAND3X1 NAND3X1_3223 ( .gnd(gnd), .vdd(vdd), .A(_13740_), .B(_14232_), .C(_14237_), .Y(_14245_) );
NAND3X1 NAND3X1_3224 ( .gnd(gnd), .vdd(vdd), .A(_13746_), .B(_14240_), .C(_14239_), .Y(_14246_) );
AOI21X1 AOI21X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_14245_), .B(_14246_), .C(_14244_), .Y(_14247_) );
INVX1 INVX1_1999 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_154_), .Y(_14248_) );
NAND2X1 NAND2X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_14248_), .B(_14223_), .Y(_14249_) );
NOR2X1 NOR2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_14248_), .B(_14223_), .Y(_14250_) );
INVX2 INVX2_504 ( .gnd(gnd), .vdd(vdd), .A(_14250_), .Y(_14251_) );
NAND3X1 NAND3X1_3225 ( .gnd(gnd), .vdd(vdd), .A(_13460_), .B(_14249_), .C(_14251_), .Y(_14252_) );
INVX1 INVX1_2000 ( .gnd(gnd), .vdd(vdd), .A(_14249_), .Y(_14253_) );
OAI21X1 OAI21X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_14253_), .B(_14250_), .C(_13461_), .Y(_14254_) );
NAND3X1 NAND3X1_3226 ( .gnd(gnd), .vdd(vdd), .A(_13464_), .B(_14254_), .C(_14252_), .Y(_14255_) );
NAND2X1 NAND2X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_14254_), .B(_14252_), .Y(_14256_) );
OAI21X1 OAI21X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_13388_), .B(_13462_), .C(_14256_), .Y(_14257_) );
NAND2X1 NAND2X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_14255_), .B(_14257_), .Y(_14258_) );
INVX1 INVX1_2001 ( .gnd(gnd), .vdd(vdd), .A(_14258_), .Y(_14259_) );
OAI21X1 OAI21X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_14242_), .B(_14247_), .C(_14259_), .Y(_14260_) );
NAND3X1 NAND3X1_3227 ( .gnd(gnd), .vdd(vdd), .A(_14244_), .B(_14245_), .C(_14246_), .Y(_14261_) );
AOI21X1 AOI21X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_14240_), .B(_14239_), .C(_13746_), .Y(_14262_) );
AOI21X1 AOI21X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_14232_), .B(_14237_), .C(_13740_), .Y(_14263_) );
OAI21X1 OAI21X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_14262_), .B(_14263_), .C(_13873_), .Y(_14264_) );
NAND3X1 NAND3X1_3228 ( .gnd(gnd), .vdd(vdd), .A(_14258_), .B(_14261_), .C(_14264_), .Y(_14265_) );
NAND3X1 NAND3X1_3229 ( .gnd(gnd), .vdd(vdd), .A(_13871_), .B(_14265_), .C(_14260_), .Y(_14266_) );
NAND2X1 NAND2X1_1872 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_182_), .B(_14266_), .Y(_14267_) );
INVX2 INVX2_505 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_182_), .Y(_14268_) );
NAND3X1 NAND3X1_3230 ( .gnd(gnd), .vdd(vdd), .A(_14259_), .B(_14261_), .C(_14264_), .Y(_14269_) );
OAI21X1 OAI21X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_14242_), .B(_14247_), .C(_14258_), .Y(_14270_) );
AOI21X1 AOI21X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_14269_), .B(_14270_), .C(_16499_), .Y(_14271_) );
NAND2X1 NAND2X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_14268_), .B(_14271_), .Y(_14272_) );
NAND3X1 NAND3X1_3231 ( .gnd(gnd), .vdd(vdd), .A(_13757_), .B(_14267_), .C(_14272_), .Y(_14273_) );
NAND2X1 NAND2X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_14269_), .B(_14270_), .Y(_14274_) );
NAND3X1 NAND3X1_3232 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_182_), .B(_13871_), .C(_14274_), .Y(_14275_) );
NAND2X1 NAND2X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_14268_), .B(_14266_), .Y(_14276_) );
NAND3X1 NAND3X1_3233 ( .gnd(gnd), .vdd(vdd), .A(_13764_), .B(_14275_), .C(_14276_), .Y(_14277_) );
NAND3X1 NAND3X1_3234 ( .gnd(gnd), .vdd(vdd), .A(_14277_), .B(_13870_), .C(_14273_), .Y(_14278_) );
AOI21X1 AOI21X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_13757_), .B(_13762_), .C(_13267_), .Y(_14279_) );
AOI21X1 AOI21X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_13770_), .B(_13768_), .C(_14279_), .Y(_14280_) );
AOI21X1 AOI21X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_14275_), .B(_14276_), .C(_13764_), .Y(_14281_) );
AOI21X1 AOI21X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_14267_), .B(_14272_), .C(_13757_), .Y(_14282_) );
OAI21X1 OAI21X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_14282_), .B(_14281_), .C(_14280_), .Y(_14283_) );
INVX1 INVX1_2002 ( .gnd(gnd), .vdd(vdd), .A(_13473_), .Y(_14284_) );
INVX1 INVX1_2003 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_170_), .Y(_14285_) );
NAND2X1 NAND2X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_14285_), .B(_14258_), .Y(_14286_) );
INVX1 INVX1_2004 ( .gnd(gnd), .vdd(vdd), .A(_14286_), .Y(_14287_) );
NOR2X1 NOR2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_14285_), .B(_14258_), .Y(_14288_) );
NOR2X1 NOR2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_14288_), .B(_14287_), .Y(_14289_) );
AND2X2 AND2X2_319 ( .gnd(gnd), .vdd(vdd), .A(_14289_), .B(_13470_), .Y(_14290_) );
OAI21X1 OAI21X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_14287_), .B(_14288_), .C(_13469_), .Y(_14291_) );
INVX1 INVX1_2005 ( .gnd(gnd), .vdd(vdd), .A(_14291_), .Y(_14292_) );
NOR2X1 NOR2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_14292_), .B(_14290_), .Y(_14293_) );
NAND2X1 NAND2X1_1877 ( .gnd(gnd), .vdd(vdd), .A(_14284_), .B(_14293_), .Y(_14294_) );
OAI21X1 OAI21X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_14290_), .B(_14292_), .C(_13473_), .Y(_14295_) );
NAND2X1 NAND2X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_14295_), .B(_14294_), .Y(_14296_) );
NAND3X1 NAND3X1_3235 ( .gnd(gnd), .vdd(vdd), .A(_14278_), .B(_14296_), .C(_14283_), .Y(_14297_) );
NAND3X1 NAND3X1_3236 ( .gnd(gnd), .vdd(vdd), .A(_13764_), .B(_14267_), .C(_14272_), .Y(_14298_) );
NAND3X1 NAND3X1_3237 ( .gnd(gnd), .vdd(vdd), .A(_13757_), .B(_14275_), .C(_14276_), .Y(_14299_) );
AOI21X1 AOI21X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_14299_), .B(_14298_), .C(_14280_), .Y(_14300_) );
AOI21X1 AOI21X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_14277_), .B(_14273_), .C(_13870_), .Y(_14301_) );
INVX1 INVX1_2006 ( .gnd(gnd), .vdd(vdd), .A(_14296_), .Y(_14302_) );
OAI21X1 OAI21X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_14300_), .B(_14301_), .C(_14302_), .Y(_14303_) );
NAND3X1 NAND3X1_3238 ( .gnd(gnd), .vdd(vdd), .A(_13868_), .B(_14297_), .C(_14303_), .Y(_14304_) );
NAND2X1 NAND2X1_1879 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_198_), .B(_14304_), .Y(_14305_) );
INVX2 INVX2_506 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_198_), .Y(_14306_) );
AOI21X1 AOI21X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_14278_), .B(_14283_), .C(_14296_), .Y(_14307_) );
NOR2X1 NOR2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_13867_), .B(_14307_), .Y(_14308_) );
NAND3X1 NAND3X1_3239 ( .gnd(gnd), .vdd(vdd), .A(_14306_), .B(_14297_), .C(_14308_), .Y(_14309_) );
NAND3X1 NAND3X1_3240 ( .gnd(gnd), .vdd(vdd), .A(_13783_), .B(_14305_), .C(_14309_), .Y(_14310_) );
NAND3X1 NAND3X1_3241 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_198_), .B(_14297_), .C(_14308_), .Y(_14311_) );
NAND2X1 NAND2X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_14306_), .B(_14304_), .Y(_14312_) );
NAND3X1 NAND3X1_3242 ( .gnd(gnd), .vdd(vdd), .A(_13777_), .B(_14312_), .C(_14311_), .Y(_14313_) );
AOI21X1 AOI21X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_14310_), .B(_14313_), .C(_13866_), .Y(_14314_) );
NOR3X1 NOR3X1_418 ( .gnd(gnd), .vdd(vdd), .A(_13784_), .B(_13516_), .C(_13783_), .Y(_14315_) );
OAI21X1 OAI21X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_14315_), .B(_13515_), .C(_13788_), .Y(_14316_) );
NAND3X1 NAND3X1_3243 ( .gnd(gnd), .vdd(vdd), .A(_13777_), .B(_14305_), .C(_14309_), .Y(_14317_) );
NAND3X1 NAND3X1_3244 ( .gnd(gnd), .vdd(vdd), .A(_13783_), .B(_14312_), .C(_14311_), .Y(_14318_) );
AOI21X1 AOI21X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_14317_), .B(_14318_), .C(_14316_), .Y(_14319_) );
INVX1 INVX1_2007 ( .gnd(gnd), .vdd(vdd), .A(_13481_), .Y(_14320_) );
INVX1 INVX1_2008 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_186_), .Y(_14321_) );
NAND2X1 NAND2X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_14321_), .B(_14296_), .Y(_14322_) );
NOR2X1 NOR2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_14321_), .B(_14296_), .Y(_14323_) );
INVX1 INVX1_2009 ( .gnd(gnd), .vdd(vdd), .A(_14323_), .Y(_14324_) );
NAND3X1 NAND3X1_3245 ( .gnd(gnd), .vdd(vdd), .A(_13478_), .B(_14322_), .C(_14324_), .Y(_14325_) );
INVX1 INVX1_2010 ( .gnd(gnd), .vdd(vdd), .A(_14322_), .Y(_14326_) );
OAI21X1 OAI21X1_2252 ( .gnd(gnd), .vdd(vdd), .A(_14326_), .B(_14323_), .C(_13477_), .Y(_14327_) );
NAND3X1 NAND3X1_3246 ( .gnd(gnd), .vdd(vdd), .A(_14320_), .B(_14327_), .C(_14325_), .Y(_14328_) );
INVX1 INVX1_2011 ( .gnd(gnd), .vdd(vdd), .A(_14325_), .Y(_14329_) );
INVX1 INVX1_2012 ( .gnd(gnd), .vdd(vdd), .A(_14327_), .Y(_14330_) );
OAI21X1 OAI21X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_14329_), .B(_14330_), .C(_13481_), .Y(_14331_) );
NAND2X1 NAND2X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_14328_), .B(_14331_), .Y(_14332_) );
INVX1 INVX1_2013 ( .gnd(gnd), .vdd(vdd), .A(_14332_), .Y(_14333_) );
OAI21X1 OAI21X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_14314_), .B(_14319_), .C(_14333_), .Y(_14334_) );
NAND3X1 NAND3X1_3247 ( .gnd(gnd), .vdd(vdd), .A(_14317_), .B(_14318_), .C(_14316_), .Y(_14335_) );
AOI21X1 AOI21X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_14312_), .B(_14311_), .C(_13783_), .Y(_14336_) );
AOI21X1 AOI21X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_14305_), .B(_14309_), .C(_13777_), .Y(_14337_) );
OAI21X1 OAI21X1_2255 ( .gnd(gnd), .vdd(vdd), .A(_14336_), .B(_14337_), .C(_13866_), .Y(_14338_) );
NAND3X1 NAND3X1_3248 ( .gnd(gnd), .vdd(vdd), .A(_14335_), .B(_14332_), .C(_14338_), .Y(_14339_) );
NAND3X1 NAND3X1_3249 ( .gnd(gnd), .vdd(vdd), .A(_13864_), .B(_14339_), .C(_14334_), .Y(_14340_) );
NAND2X1 NAND2X1_1883 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_214_), .B(_14340_), .Y(_14341_) );
INVX2 INVX2_507 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_214_), .Y(_14342_) );
OAI21X1 OAI21X1_2256 ( .gnd(gnd), .vdd(vdd), .A(_14314_), .B(_14319_), .C(_14332_), .Y(_14343_) );
NAND3X1 NAND3X1_3250 ( .gnd(gnd), .vdd(vdd), .A(_14335_), .B(_14333_), .C(_14338_), .Y(_14344_) );
AOI21X1 AOI21X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_14344_), .B(_14343_), .C(_16517_), .Y(_14345_) );
NAND2X1 NAND2X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_14342_), .B(_14345_), .Y(_14346_) );
NAND3X1 NAND3X1_3251 ( .gnd(gnd), .vdd(vdd), .A(_13802_), .B(_14341_), .C(_14346_), .Y(_14347_) );
NAND2X1 NAND2X1_1885 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_214_), .B(_14345_), .Y(_14348_) );
NAND2X1 NAND2X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_14342_), .B(_14340_), .Y(_14349_) );
NAND3X1 NAND3X1_3252 ( .gnd(gnd), .vdd(vdd), .A(_13796_), .B(_14349_), .C(_14348_), .Y(_14350_) );
AOI21X1 AOI21X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_14347_), .B(_14350_), .C(_13863_), .Y(_14351_) );
NOR3X1 NOR3X1_419 ( .gnd(gnd), .vdd(vdd), .A(_13803_), .B(_13513_), .C(_13802_), .Y(_14352_) );
OAI21X1 OAI21X1_2257 ( .gnd(gnd), .vdd(vdd), .A(_14352_), .B(_13512_), .C(_13807_), .Y(_14353_) );
NAND3X1 NAND3X1_3253 ( .gnd(gnd), .vdd(vdd), .A(_13796_), .B(_14341_), .C(_14346_), .Y(_14354_) );
NAND3X1 NAND3X1_3254 ( .gnd(gnd), .vdd(vdd), .A(_13802_), .B(_14349_), .C(_14348_), .Y(_14355_) );
AOI21X1 AOI21X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_14354_), .B(_14355_), .C(_14353_), .Y(_14356_) );
INVX1 INVX1_2014 ( .gnd(gnd), .vdd(vdd), .A(_13489_), .Y(_14357_) );
INVX1 INVX1_2015 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_202_), .Y(_14358_) );
NAND2X1 NAND2X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_14358_), .B(_14332_), .Y(_14359_) );
NOR2X1 NOR2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_14358_), .B(_14332_), .Y(_14360_) );
INVX2 INVX2_508 ( .gnd(gnd), .vdd(vdd), .A(_14360_), .Y(_14361_) );
NAND3X1 NAND3X1_3255 ( .gnd(gnd), .vdd(vdd), .A(_13486_), .B(_14359_), .C(_14361_), .Y(_14362_) );
INVX1 INVX1_2016 ( .gnd(gnd), .vdd(vdd), .A(_14359_), .Y(_14363_) );
OAI21X1 OAI21X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_14363_), .B(_14360_), .C(_13485_), .Y(_14364_) );
NAND3X1 NAND3X1_3256 ( .gnd(gnd), .vdd(vdd), .A(_14357_), .B(_14364_), .C(_14362_), .Y(_14365_) );
INVX1 INVX1_2017 ( .gnd(gnd), .vdd(vdd), .A(_14362_), .Y(_14366_) );
INVX1 INVX1_2018 ( .gnd(gnd), .vdd(vdd), .A(_14364_), .Y(_14367_) );
OAI21X1 OAI21X1_2259 ( .gnd(gnd), .vdd(vdd), .A(_14366_), .B(_14367_), .C(_13489_), .Y(_14368_) );
NAND2X1 NAND2X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_14365_), .B(_14368_), .Y(_14369_) );
INVX2 INVX2_509 ( .gnd(gnd), .vdd(vdd), .A(_14369_), .Y(_14370_) );
OAI21X1 OAI21X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_14356_), .B(_14351_), .C(_14370_), .Y(_14371_) );
NAND3X1 NAND3X1_3257 ( .gnd(gnd), .vdd(vdd), .A(_14354_), .B(_14355_), .C(_14353_), .Y(_14372_) );
AOI21X1 AOI21X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_14349_), .B(_14348_), .C(_13802_), .Y(_14373_) );
AOI21X1 AOI21X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_14341_), .B(_14346_), .C(_13796_), .Y(_14374_) );
OAI21X1 OAI21X1_2261 ( .gnd(gnd), .vdd(vdd), .A(_14373_), .B(_14374_), .C(_13863_), .Y(_14375_) );
NAND3X1 NAND3X1_3258 ( .gnd(gnd), .vdd(vdd), .A(_14369_), .B(_14375_), .C(_14372_), .Y(_14376_) );
NAND3X1 NAND3X1_3259 ( .gnd(gnd), .vdd(vdd), .A(_13861_), .B(_14376_), .C(_14371_), .Y(_14377_) );
NAND2X1 NAND2X1_1889 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_230_), .B(_14377_), .Y(_14378_) );
INVX2 INVX2_510 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_230_), .Y(_14379_) );
OAI21X1 OAI21X1_2262 ( .gnd(gnd), .vdd(vdd), .A(_14356_), .B(_14351_), .C(_14369_), .Y(_14380_) );
NAND3X1 NAND3X1_3260 ( .gnd(gnd), .vdd(vdd), .A(_14370_), .B(_14375_), .C(_14372_), .Y(_14381_) );
AOI21X1 AOI21X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_14381_), .B(_14380_), .C(_13860_), .Y(_14382_) );
NAND2X1 NAND2X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_14379_), .B(_14382_), .Y(_14383_) );
NAND3X1 NAND3X1_3261 ( .gnd(gnd), .vdd(vdd), .A(_13821_), .B(_14378_), .C(_14383_), .Y(_14384_) );
NAND2X1 NAND2X1_1891 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_230_), .B(_14382_), .Y(_14385_) );
NAND2X1 NAND2X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_14379_), .B(_14377_), .Y(_14386_) );
NAND3X1 NAND3X1_3262 ( .gnd(gnd), .vdd(vdd), .A(_13815_), .B(_14386_), .C(_14385_), .Y(_14387_) );
AOI21X1 AOI21X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_14384_), .B(_14387_), .C(_13857_), .Y(_14388_) );
NOR3X1 NOR3X1_420 ( .gnd(gnd), .vdd(vdd), .A(_13822_), .B(_13510_), .C(_13821_), .Y(_14389_) );
OAI21X1 OAI21X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_14389_), .B(_13509_), .C(_13826_), .Y(_14390_) );
NAND3X1 NAND3X1_3263 ( .gnd(gnd), .vdd(vdd), .A(_13815_), .B(_14378_), .C(_14383_), .Y(_14391_) );
NAND3X1 NAND3X1_3264 ( .gnd(gnd), .vdd(vdd), .A(_13821_), .B(_14386_), .C(_14385_), .Y(_14392_) );
AOI21X1 AOI21X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_14391_), .B(_14392_), .C(_14390_), .Y(_14393_) );
INVX1 INVX1_2019 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .Y(_14394_) );
INVX1 INVX1_2020 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_218_), .Y(_14395_) );
NAND2X1 NAND2X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_14395_), .B(_14369_), .Y(_14396_) );
NOR2X1 NOR2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_14395_), .B(_14369_), .Y(_14397_) );
INVX2 INVX2_511 ( .gnd(gnd), .vdd(vdd), .A(_14397_), .Y(_14398_) );
NAND2X1 NAND2X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_14396_), .B(_14398_), .Y(_14399_) );
OR2X2 OR2X2_345 ( .gnd(gnd), .vdd(vdd), .A(_14399_), .B(_13493_), .Y(_14400_) );
AOI21X1 AOI21X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_14396_), .B(_14398_), .C(_13494_), .Y(_14401_) );
INVX1 INVX1_2021 ( .gnd(gnd), .vdd(vdd), .A(_14401_), .Y(_14402_) );
NAND3X1 NAND3X1_3265 ( .gnd(gnd), .vdd(vdd), .A(_14394_), .B(_14402_), .C(_14400_), .Y(_14403_) );
NOR2X1 NOR2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_13493_), .B(_14399_), .Y(_14404_) );
OAI21X1 OAI21X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_14404_), .B(_14401_), .C(_13497_), .Y(_14405_) );
NAND2X1 NAND2X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_14405_), .B(_14403_), .Y(_14406_) );
INVX2 INVX2_512 ( .gnd(gnd), .vdd(vdd), .A(_14406_), .Y(_14407_) );
OAI21X1 OAI21X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_14393_), .B(_14388_), .C(_14407_), .Y(_14408_) );
NAND3X1 NAND3X1_3266 ( .gnd(gnd), .vdd(vdd), .A(_14391_), .B(_14392_), .C(_14390_), .Y(_14409_) );
AOI21X1 AOI21X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_14386_), .B(_14385_), .C(_13821_), .Y(_14410_) );
AOI21X1 AOI21X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_14378_), .B(_14383_), .C(_13815_), .Y(_14411_) );
OAI21X1 OAI21X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_14410_), .B(_14411_), .C(_13857_), .Y(_14412_) );
NAND3X1 NAND3X1_3267 ( .gnd(gnd), .vdd(vdd), .A(_14412_), .B(_14406_), .C(_14409_), .Y(_14413_) );
NAND3X1 NAND3X1_3268 ( .gnd(gnd), .vdd(vdd), .A(_16767_), .B(_14413_), .C(_14408_), .Y(_14414_) );
NAND2X1 NAND2X1_1896 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_246_), .B(_14414_), .Y(_14415_) );
INVX1 INVX1_2022 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_246_), .Y(_14416_) );
NAND3X1 NAND3X1_3269 ( .gnd(gnd), .vdd(vdd), .A(_14412_), .B(_14407_), .C(_14409_), .Y(_14417_) );
OAI21X1 OAI21X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_14393_), .B(_14388_), .C(_14406_), .Y(_14418_) );
AOI21X1 AOI21X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_14417_), .B(_14418_), .C(_16539_), .Y(_14419_) );
NAND2X1 NAND2X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_14416_), .B(_14419_), .Y(_14420_) );
NAND3X1 NAND3X1_3270 ( .gnd(gnd), .vdd(vdd), .A(_13840_), .B(_14415_), .C(_14420_), .Y(_14421_) );
NAND2X1 NAND2X1_1898 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_246_), .B(_14419_), .Y(_14422_) );
NAND2X1 NAND2X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_14416_), .B(_14414_), .Y(_14423_) );
NAND3X1 NAND3X1_3271 ( .gnd(gnd), .vdd(vdd), .A(_13832_), .B(_14423_), .C(_14422_), .Y(_14424_) );
AOI21X1 AOI21X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_14421_), .B(_14424_), .C(_13855_), .Y(_14425_) );
OAI21X1 OAI21X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_13845_), .B(_13844_), .C(_13842_), .Y(_14426_) );
NAND3X1 NAND3X1_3272 ( .gnd(gnd), .vdd(vdd), .A(_13832_), .B(_14415_), .C(_14420_), .Y(_14427_) );
NAND3X1 NAND3X1_3273 ( .gnd(gnd), .vdd(vdd), .A(_13840_), .B(_14423_), .C(_14422_), .Y(_14428_) );
AOI21X1 AOI21X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_14427_), .B(_14428_), .C(_14426_), .Y(_14429_) );
INVX1 INVX1_2023 ( .gnd(gnd), .vdd(vdd), .A(_13505_), .Y(_14430_) );
NOR2X1 NOR2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_234_), .B(_14407_), .Y(_14431_) );
INVX1 INVX1_2024 ( .gnd(gnd), .vdd(vdd), .A(_14431_), .Y(_14432_) );
NAND2X1 NAND2X1_1900 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_234_), .B(_14407_), .Y(_14433_) );
NAND3X1 NAND3X1_3274 ( .gnd(gnd), .vdd(vdd), .A(_13502_), .B(_14433_), .C(_14432_), .Y(_14434_) );
INVX2 INVX2_513 ( .gnd(gnd), .vdd(vdd), .A(_14433_), .Y(_14435_) );
OAI21X1 OAI21X1_2269 ( .gnd(gnd), .vdd(vdd), .A(_14435_), .B(_14431_), .C(_13501_), .Y(_14436_) );
NAND3X1 NAND3X1_3275 ( .gnd(gnd), .vdd(vdd), .A(_14430_), .B(_14436_), .C(_14434_), .Y(_14437_) );
NOR3X1 NOR3X1_421 ( .gnd(gnd), .vdd(vdd), .A(_13501_), .B(_14431_), .C(_14435_), .Y(_14438_) );
AOI21X1 AOI21X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_14433_), .B(_14432_), .C(_13502_), .Y(_14439_) );
OAI21X1 OAI21X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_14439_), .B(_14438_), .C(_13505_), .Y(_14440_) );
NAND2X1 NAND2X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_14437_), .B(_14440_), .Y(_14441_) );
INVX2 INVX2_514 ( .gnd(gnd), .vdd(vdd), .A(_14441_), .Y(_14442_) );
OAI21X1 OAI21X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_14429_), .B(_14425_), .C(_14442_), .Y(_14443_) );
NAND3X1 NAND3X1_3276 ( .gnd(gnd), .vdd(vdd), .A(_14427_), .B(_14428_), .C(_14426_), .Y(_14444_) );
NAND3X1 NAND3X1_3277 ( .gnd(gnd), .vdd(vdd), .A(_14421_), .B(_14424_), .C(_13855_), .Y(_14445_) );
NAND3X1 NAND3X1_3278 ( .gnd(gnd), .vdd(vdd), .A(_14445_), .B(_14441_), .C(_14444_), .Y(_14446_) );
NAND2X1 NAND2X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_14446_), .B(_14443_), .Y(_14447_) );
XOR2X1 XOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_14447_), .B(_13854_), .Y(module_3_H_6_) );
OAI21X1 OAI21X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_14429_), .B(_14425_), .C(_14441_), .Y(_14448_) );
NAND3X1 NAND3X1_3279 ( .gnd(gnd), .vdd(vdd), .A(_14445_), .B(_14442_), .C(_14444_), .Y(_14449_) );
NAND3X1 NAND3X1_3280 ( .gnd(gnd), .vdd(vdd), .A(_14449_), .B(_14448_), .C(_13854_), .Y(_14450_) );
AOI21X1 AOI21X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_14423_), .B(_14422_), .C(_13840_), .Y(_14451_) );
AOI21X1 AOI21X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_14428_), .B(_14426_), .C(_14451_), .Y(_14452_) );
AOI21X1 AOI21X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_14430_), .B(_14436_), .C(_14438_), .Y(_14453_) );
OAI21X1 OAI21X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(_14401_), .C(_14400_), .Y(_14454_) );
AOI21X1 AOI21X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_14357_), .B(_14364_), .C(_14366_), .Y(_14455_) );
INVX1 INVX1_2025 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_203_), .Y(_14456_) );
OAI21X1 OAI21X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_14330_), .B(_13481_), .C(_14325_), .Y(_14457_) );
INVX1 INVX1_2026 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_187_), .Y(_14458_) );
AOI21X1 AOI21X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_14284_), .B(_14291_), .C(_14290_), .Y(_14459_) );
INVX1 INVX1_2027 ( .gnd(gnd), .vdd(vdd), .A(_14459_), .Y(_14460_) );
INVX1 INVX1_2028 ( .gnd(gnd), .vdd(vdd), .A(_14288_), .Y(_14461_) );
INVX1 INVX1_2029 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_171_), .Y(_14462_) );
OAI21X1 OAI21X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_14256_), .B(_13465_), .C(_14252_), .Y(_14463_) );
INVX1 INVX1_2030 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_155_), .Y(_14464_) );
AOI21X1 AOI21X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_13456_), .B(_14219_), .C(_14217_), .Y(_14465_) );
INVX1 INVX1_2031 ( .gnd(gnd), .vdd(vdd), .A(_14183_), .Y(_14466_) );
OAI21X1 OAI21X1_2276 ( .gnd(gnd), .vdd(vdd), .A(_14466_), .B(_13449_), .C(_14180_), .Y(_14467_) );
OAI21X1 OAI21X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_13442_), .B(_14142_), .C(_14145_), .Y(_14468_) );
INVX1 INVX1_2032 ( .gnd(gnd), .vdd(vdd), .A(_14138_), .Y(_14469_) );
OAI21X1 OAI21X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_13436_), .B(_14102_), .C(_14105_), .Y(_14470_) );
AOI21X1 AOI21X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_14063_), .B(_14065_), .C(_14058_), .Y(_14471_) );
INVX1 INVX1_2033 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf0_), .Y(_14472_) );
NOR2X1 NOR2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .B(_13419_), .Y(_14473_) );
AOI21X1 AOI21X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_14473_), .B(_14022_), .C(_14025_), .Y(_14474_) );
INVX1 INVX1_2034 ( .gnd(gnd), .vdd(vdd), .A(_13986_), .Y(_14475_) );
AOI21X1 AOI21X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_13979_), .B(_14475_), .C(_13985_), .Y(_14476_) );
INVX1 INVX1_2035 ( .gnd(gnd), .vdd(vdd), .A(_13983_), .Y(_14477_) );
INVX1 INVX1_2036 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .Y(_14478_) );
OAI21X1 OAI21X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_13953_), .B(_13950_), .C(_13946_), .Y(_14479_) );
NOR2X1 NOR2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_27_), .B(module_3_W_11_), .Y(_14480_) );
INVX1 INVX1_2037 ( .gnd(gnd), .vdd(vdd), .A(_14480_), .Y(_14481_) );
NAND2X1 NAND2X1_1903 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_27_), .B(module_3_W_11_), .Y(_14482_) );
NAND2X1 NAND2X1_1904 ( .gnd(gnd), .vdd(vdd), .A(_14482_), .B(_14481_), .Y(_14483_) );
NAND3X1 NAND3X1_3281 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_26_), .B(module_3_W_10_), .C(_14483_), .Y(_14484_) );
NAND3X1 NAND3X1_3282 ( .gnd(gnd), .vdd(vdd), .A(_13942_), .B(_14482_), .C(_14481_), .Y(_14485_) );
NAND2X1 NAND2X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_14485_), .B(_14484_), .Y(_14486_) );
XOR2X1 XOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_14479_), .B(_14486_), .Y(_14487_) );
NAND2X1 NAND2X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_14478_), .B(_14487_), .Y(_14488_) );
XNOR2X1 XNOR2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_14479_), .B(_14486_), .Y(_14489_) );
NAND2X1 NAND2X1_1907 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .B(_14489_), .Y(_14490_) );
NAND2X1 NAND2X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_14490_), .B(_14488_), .Y(_14491_) );
NAND2X1 NAND2X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_14477_), .B(_14491_), .Y(_14492_) );
NAND3X1 NAND3X1_3283 ( .gnd(gnd), .vdd(vdd), .A(_13983_), .B(_14490_), .C(_14488_), .Y(_14493_) );
NAND2X1 NAND2X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_14493_), .B(_14492_), .Y(_14494_) );
XNOR2X1 XNOR2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_14494_), .B(_14476_), .Y(_14495_) );
NAND2X1 NAND2X1_1911 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf3_), .B(_14495_), .Y(_14496_) );
INVX1 INVX1_2038 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf2_), .Y(_14497_) );
OR2X2 OR2X2_346 ( .gnd(gnd), .vdd(vdd), .A(_13984_), .B(_13980_), .Y(_14498_) );
OAI21X1 OAI21X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_13414_), .B(_13986_), .C(_14498_), .Y(_14499_) );
XNOR2X1 XNOR2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_14494_), .B(_14499_), .Y(_14500_) );
NAND2X1 NAND2X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_14497_), .B(_14500_), .Y(_14501_) );
NAND2X1 NAND2X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_14496_), .B(_14501_), .Y(_14502_) );
NOR2X1 NOR2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_14017_), .B(_14502_), .Y(_14503_) );
AOI21X1 AOI21X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_14496_), .B(_14501_), .C(_14021_), .Y(_14504_) );
OAI21X1 OAI21X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_14503_), .B(_14504_), .C(_14474_), .Y(_14505_) );
OAI21X1 OAI21X1_2282 ( .gnd(gnd), .vdd(vdd), .A(_14026_), .B(_13420_), .C(_14018_), .Y(_14506_) );
OR2X2 OR2X2_347 ( .gnd(gnd), .vdd(vdd), .A(_14502_), .B(_14017_), .Y(_14507_) );
INVX1 INVX1_2039 ( .gnd(gnd), .vdd(vdd), .A(_14504_), .Y(_14508_) );
NAND3X1 NAND3X1_3284 ( .gnd(gnd), .vdd(vdd), .A(_14508_), .B(_14506_), .C(_14507_), .Y(_14509_) );
NAND2X1 NAND2X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_14505_), .B(_14509_), .Y(_14510_) );
NAND2X1 NAND2X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_14472_), .B(_14510_), .Y(_14511_) );
AND2X2 AND2X2_320 ( .gnd(gnd), .vdd(vdd), .A(_14509_), .B(_14505_), .Y(_14512_) );
NAND2X1 NAND2X1_1916 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf3_), .B(_14512_), .Y(_14513_) );
AOI21X1 AOI21X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_14511_), .B(_14513_), .C(_14060_), .Y(_14514_) );
NAND3X1 NAND3X1_3285 ( .gnd(gnd), .vdd(vdd), .A(_14060_), .B(_14511_), .C(_14513_), .Y(_14515_) );
INVX2 INVX2_515 ( .gnd(gnd), .vdd(vdd), .A(_14515_), .Y(_14516_) );
OAI21X1 OAI21X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_14516_), .B(_14514_), .C(_14471_), .Y(_14517_) );
INVX2 INVX2_516 ( .gnd(gnd), .vdd(vdd), .A(_14517_), .Y(_14518_) );
NOR2X1 NOR2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_14514_), .B(_14516_), .Y(_14519_) );
OAI21X1 OAI21X1_2284 ( .gnd(gnd), .vdd(vdd), .A(_14058_), .B(_14062_), .C(_14519_), .Y(_14520_) );
INVX2 INVX2_517 ( .gnd(gnd), .vdd(vdd), .A(_14520_), .Y(_14521_) );
OAI21X1 OAI21X1_2285 ( .gnd(gnd), .vdd(vdd), .A(_14521_), .B(_14518_), .C(bloque_datos_59_bF_buf1_), .Y(_14522_) );
INVX1 INVX1_2040 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf0_), .Y(_14523_) );
NAND3X1 NAND3X1_3286 ( .gnd(gnd), .vdd(vdd), .A(_14523_), .B(_14517_), .C(_14520_), .Y(_14524_) );
NAND3X1 NAND3X1_3287 ( .gnd(gnd), .vdd(vdd), .A(_14098_), .B(_14524_), .C(_14522_), .Y(_14525_) );
OAI21X1 OAI21X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_14521_), .B(_14518_), .C(_14523_), .Y(_14526_) );
NAND3X1 NAND3X1_3288 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf4_), .B(_14517_), .C(_14520_), .Y(_14527_) );
NAND3X1 NAND3X1_3289 ( .gnd(gnd), .vdd(vdd), .A(_14101_), .B(_14527_), .C(_14526_), .Y(_14528_) );
AOI21X1 AOI21X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_14525_), .B(_14528_), .C(_14470_), .Y(_14529_) );
NAND3X1 NAND3X1_3290 ( .gnd(gnd), .vdd(vdd), .A(_14470_), .B(_14525_), .C(_14528_), .Y(_14530_) );
INVX2 INVX2_518 ( .gnd(gnd), .vdd(vdd), .A(_14530_), .Y(_14531_) );
OAI21X1 OAI21X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_14531_), .B(_14529_), .C(bloque_datos_75_bF_buf3_), .Y(_14532_) );
INVX1 INVX1_2041 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf2_), .Y(_14533_) );
INVX1 INVX1_2042 ( .gnd(gnd), .vdd(vdd), .A(_14529_), .Y(_14534_) );
NAND3X1 NAND3X1_3291 ( .gnd(gnd), .vdd(vdd), .A(_14533_), .B(_14530_), .C(_14534_), .Y(_14535_) );
NAND3X1 NAND3X1_3292 ( .gnd(gnd), .vdd(vdd), .A(_14469_), .B(_14535_), .C(_14532_), .Y(_14536_) );
OAI21X1 OAI21X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_14531_), .B(_14529_), .C(_14533_), .Y(_14537_) );
NAND3X1 NAND3X1_3293 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf1_), .B(_14530_), .C(_14534_), .Y(_14538_) );
NAND3X1 NAND3X1_3294 ( .gnd(gnd), .vdd(vdd), .A(_14138_), .B(_14538_), .C(_14537_), .Y(_14539_) );
AOI21X1 AOI21X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_14536_), .B(_14539_), .C(_14468_), .Y(_14540_) );
NAND3X1 NAND3X1_3295 ( .gnd(gnd), .vdd(vdd), .A(_14468_), .B(_14536_), .C(_14539_), .Y(_14541_) );
INVX2 INVX2_519 ( .gnd(gnd), .vdd(vdd), .A(_14541_), .Y(_14542_) );
OAI21X1 OAI21X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_14542_), .B(_14540_), .C(bloque_datos_91_bF_buf0_), .Y(_14543_) );
INVX1 INVX1_2043 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf3_), .Y(_14544_) );
INVX1 INVX1_2044 ( .gnd(gnd), .vdd(vdd), .A(_14540_), .Y(_14545_) );
NAND3X1 NAND3X1_3296 ( .gnd(gnd), .vdd(vdd), .A(_14544_), .B(_14541_), .C(_14545_), .Y(_14546_) );
NAND3X1 NAND3X1_3297 ( .gnd(gnd), .vdd(vdd), .A(_14182_), .B(_14546_), .C(_14543_), .Y(_14547_) );
OAI21X1 OAI21X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_14542_), .B(_14540_), .C(_14544_), .Y(_14548_) );
NAND3X1 NAND3X1_3298 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf2_), .B(_14541_), .C(_14545_), .Y(_14549_) );
NAND3X1 NAND3X1_3299 ( .gnd(gnd), .vdd(vdd), .A(_14179_), .B(_14549_), .C(_14548_), .Y(_14550_) );
NAND3X1 NAND3X1_3300 ( .gnd(gnd), .vdd(vdd), .A(_14547_), .B(_14550_), .C(_14467_), .Y(_14551_) );
INVX1 INVX1_2045 ( .gnd(gnd), .vdd(vdd), .A(_14551_), .Y(_14552_) );
AOI21X1 AOI21X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_14547_), .B(_14550_), .C(_14467_), .Y(_14553_) );
NOR2X1 NOR2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_14553_), .B(_14552_), .Y(_14554_) );
XNOR2X1 XNOR2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_14554_), .B(module_3_W_139_), .Y(_14555_) );
NOR2X1 NOR2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_14215_), .B(_14555_), .Y(_14556_) );
INVX1 INVX1_2046 ( .gnd(gnd), .vdd(vdd), .A(_14556_), .Y(_14557_) );
OAI21X1 OAI21X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_14213_), .B(_14189_), .C(_14555_), .Y(_14558_) );
NAND2X1 NAND2X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_14558_), .B(_14557_), .Y(_14559_) );
OR2X2 OR2X2_348 ( .gnd(gnd), .vdd(vdd), .A(_14559_), .B(_14465_), .Y(_14560_) );
INVX1 INVX1_2047 ( .gnd(gnd), .vdd(vdd), .A(_14558_), .Y(_14561_) );
OAI21X1 OAI21X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_14561_), .B(_14556_), .C(_14465_), .Y(_14562_) );
NAND2X1 NAND2X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_14562_), .B(_14560_), .Y(_14563_) );
NAND2X1 NAND2X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_14464_), .B(_14563_), .Y(_14564_) );
INVX1 INVX1_2048 ( .gnd(gnd), .vdd(vdd), .A(_14564_), .Y(_14565_) );
NOR2X1 NOR2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_14464_), .B(_14563_), .Y(_14566_) );
NOR3X1 NOR3X1_422 ( .gnd(gnd), .vdd(vdd), .A(_14251_), .B(_14566_), .C(_14565_), .Y(_14567_) );
INVX2 INVX2_520 ( .gnd(gnd), .vdd(vdd), .A(_14566_), .Y(_14568_) );
AOI21X1 AOI21X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_14564_), .B(_14568_), .C(_14250_), .Y(_14569_) );
NOR2X1 NOR2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_14567_), .B(_14569_), .Y(_14570_) );
AND2X2 AND2X2_321 ( .gnd(gnd), .vdd(vdd), .A(_14570_), .B(_14463_), .Y(_14571_) );
AND2X2 AND2X2_322 ( .gnd(gnd), .vdd(vdd), .A(_14255_), .B(_14252_), .Y(_14572_) );
OAI21X1 OAI21X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_14569_), .B(_14567_), .C(_14572_), .Y(_14573_) );
INVX2 INVX2_521 ( .gnd(gnd), .vdd(vdd), .A(_14573_), .Y(_14574_) );
OAI21X1 OAI21X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_14571_), .B(_14574_), .C(_14462_), .Y(_14575_) );
NOR2X1 NOR2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_14574_), .B(_14571_), .Y(_14576_) );
NAND2X1 NAND2X1_1920 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_171_), .B(_14576_), .Y(_14577_) );
NAND2X1 NAND2X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_14575_), .B(_14577_), .Y(_14578_) );
NOR2X1 NOR2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_14461_), .B(_14578_), .Y(_14579_) );
AOI21X1 AOI21X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_14575_), .B(_14577_), .C(_14288_), .Y(_14580_) );
NOR2X1 NOR2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_14580_), .B(_14579_), .Y(_14581_) );
AND2X2 AND2X2_323 ( .gnd(gnd), .vdd(vdd), .A(_14581_), .B(_14460_), .Y(_14582_) );
OAI21X1 OAI21X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_14579_), .B(_14580_), .C(_14459_), .Y(_14583_) );
INVX2 INVX2_522 ( .gnd(gnd), .vdd(vdd), .A(_14583_), .Y(_14584_) );
OAI21X1 OAI21X1_2296 ( .gnd(gnd), .vdd(vdd), .A(_14582_), .B(_14584_), .C(_14458_), .Y(_14585_) );
NOR2X1 NOR2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_14584_), .B(_14582_), .Y(_14586_) );
NAND2X1 NAND2X1_1922 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_187_), .B(_14586_), .Y(_14587_) );
NAND3X1 NAND3X1_3301 ( .gnd(gnd), .vdd(vdd), .A(_14323_), .B(_14585_), .C(_14587_), .Y(_14588_) );
INVX2 INVX2_523 ( .gnd(gnd), .vdd(vdd), .A(_14588_), .Y(_14589_) );
AOI21X1 AOI21X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_14585_), .B(_14587_), .C(_14323_), .Y(_14590_) );
NOR2X1 NOR2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_14590_), .B(_14589_), .Y(_14591_) );
NAND2X1 NAND2X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_14457_), .B(_14591_), .Y(_14592_) );
AOI21X1 AOI21X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_14320_), .B(_14327_), .C(_14329_), .Y(_14593_) );
OAI21X1 OAI21X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_14589_), .B(_14590_), .C(_14593_), .Y(_14594_) );
NAND2X1 NAND2X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_14594_), .B(_14592_), .Y(_14595_) );
NAND2X1 NAND2X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_14456_), .B(_14595_), .Y(_14596_) );
NOR2X1 NOR2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_14456_), .B(_14595_), .Y(_14597_) );
INVX2 INVX2_524 ( .gnd(gnd), .vdd(vdd), .A(_14597_), .Y(_14598_) );
NAND3X1 NAND3X1_3302 ( .gnd(gnd), .vdd(vdd), .A(_14360_), .B(_14596_), .C(_14598_), .Y(_14599_) );
INVX1 INVX1_2049 ( .gnd(gnd), .vdd(vdd), .A(_14596_), .Y(_14600_) );
OAI21X1 OAI21X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_14600_), .B(_14597_), .C(_14361_), .Y(_14601_) );
NAND2X1 NAND2X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_14601_), .B(_14599_), .Y(_14602_) );
NOR2X1 NOR2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_14455_), .B(_14602_), .Y(_14603_) );
OAI21X1 OAI21X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_14367_), .B(_13489_), .C(_14362_), .Y(_14604_) );
AOI21X1 AOI21X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_14601_), .B(_14599_), .C(_14604_), .Y(_14605_) );
NOR2X1 NOR2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_14605_), .B(_14603_), .Y(_14606_) );
NOR2X1 NOR2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_219_), .B(_14606_), .Y(_14607_) );
AND2X2 AND2X2_324 ( .gnd(gnd), .vdd(vdd), .A(_14606_), .B(module_3_W_219_), .Y(_14608_) );
NOR3X1 NOR3X1_423 ( .gnd(gnd), .vdd(vdd), .A(_14607_), .B(_14398_), .C(_14608_), .Y(_14609_) );
OR2X2 OR2X2_349 ( .gnd(gnd), .vdd(vdd), .A(_14606_), .B(module_3_W_219_), .Y(_14610_) );
NAND2X1 NAND2X1_1927 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_219_), .B(_14606_), .Y(_14611_) );
AOI21X1 AOI21X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_14611_), .B(_14610_), .C(_14397_), .Y(_14612_) );
NOR2X1 NOR2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_14612_), .B(_14609_), .Y(_14613_) );
AND2X2 AND2X2_325 ( .gnd(gnd), .vdd(vdd), .A(_14613_), .B(_14454_), .Y(_14614_) );
NOR2X1 NOR2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_14454_), .B(_14613_), .Y(_14615_) );
NOR2X1 NOR2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_14615_), .B(_14614_), .Y(_14616_) );
OR2X2 OR2X2_350 ( .gnd(gnd), .vdd(vdd), .A(_14616_), .B(module_3_W_235_), .Y(_14617_) );
NAND2X1 NAND2X1_1928 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_235_), .B(_14616_), .Y(_14618_) );
NAND3X1 NAND3X1_3303 ( .gnd(gnd), .vdd(vdd), .A(_14435_), .B(_14618_), .C(_14617_), .Y(_14619_) );
INVX2 INVX2_525 ( .gnd(gnd), .vdd(vdd), .A(_14619_), .Y(_14620_) );
AOI21X1 AOI21X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_14618_), .B(_14617_), .C(_14435_), .Y(_14621_) );
OAI21X1 OAI21X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_14620_), .B(_14621_), .C(_14453_), .Y(_14622_) );
INVX1 INVX1_2050 ( .gnd(gnd), .vdd(vdd), .A(_14622_), .Y(_14623_) );
OAI21X1 OAI21X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_14439_), .B(_13505_), .C(_14434_), .Y(_14624_) );
NOR2X1 NOR2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_14621_), .B(_14620_), .Y(_14625_) );
AND2X2 AND2X2_326 ( .gnd(gnd), .vdd(vdd), .A(_14625_), .B(_14624_), .Y(_14626_) );
NOR2X1 NOR2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_14623_), .B(_14626_), .Y(_14627_) );
INVX2 INVX2_526 ( .gnd(gnd), .vdd(vdd), .A(_14627_), .Y(_14628_) );
INVX1 INVX1_2051 ( .gnd(gnd), .vdd(vdd), .A(_14616_), .Y(_14629_) );
AOI21X1 AOI21X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_14318_), .B(_14316_), .C(_14336_), .Y(_14630_) );
OAI21X1 OAI21X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_14282_), .B(_14280_), .C(_14273_), .Y(_14631_) );
INVX1 INVX1_2052 ( .gnd(gnd), .vdd(vdd), .A(_14631_), .Y(_14632_) );
OR2X2 OR2X2_351 ( .gnd(gnd), .vdd(vdd), .A(_14582_), .B(_14584_), .Y(_14633_) );
OAI21X1 OAI21X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_14236_), .B(_14233_), .C(module_3_W_167_), .Y(_14634_) );
INVX1 INVX1_2053 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_167_), .Y(_14635_) );
NAND3X1 NAND3X1_3304 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_166_), .B(_14635_), .C(_14231_), .Y(_14636_) );
OR2X2 OR2X2_352 ( .gnd(gnd), .vdd(vdd), .A(_14571_), .B(_14574_), .Y(_14637_) );
INVX1 INVX1_2054 ( .gnd(gnd), .vdd(vdd), .A(_14160_), .Y(_14638_) );
AOI21X1 AOI21X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_13881_), .B(_14128_), .C(_14131_), .Y(_14639_) );
INVX1 INVX1_2055 ( .gnd(gnd), .vdd(vdd), .A(_14639_), .Y(_14640_) );
NOR2X1 NOR2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_14540_), .B(_14542_), .Y(_14641_) );
OAI21X1 OAI21X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_14089_), .B(_14091_), .C(_14084_), .Y(_14642_) );
NOR2X1 NOR2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_14529_), .B(_14531_), .Y(_14643_) );
OAI21X1 OAI21X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_14047_), .B(_14049_), .C(_14042_), .Y(_14644_) );
NOR2X1 NOR2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_14518_), .B(_14521_), .Y(_14645_) );
INVX1 INVX1_2056 ( .gnd(gnd), .vdd(vdd), .A(_14645_), .Y(_14646_) );
AOI21X1 AOI21X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_14007_), .B(_13887_), .C(_14010_), .Y(_14647_) );
AOI21X1 AOI21X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_13972_), .B(_13889_), .C(_13975_), .Y(_14648_) );
AOI21X1 AOI21X1_2054 ( .gnd(gnd), .vdd(vdd), .A(_13892_), .B(_13934_), .C(_13938_), .Y(_14649_) );
INVX1 INVX1_2057 ( .gnd(gnd), .vdd(vdd), .A(_13909_), .Y(_14650_) );
NOR2X1 NOR2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_14650_), .B(_13914_), .Y(_14651_) );
XNOR2X1 XNOR2X1_379 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_7_), .B(module_3_W_23_), .Y(_14652_) );
XOR2X1 XOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_16590_), .B(_14652_), .Y(_14653_) );
XNOR2X1 XNOR2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_13900_), .B(module_3_W_11_), .Y(_14654_) );
XNOR2X1 XNOR2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_14654_), .B(_14653_), .Y(_14655_) );
XNOR2X1 XNOR2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_14655_), .B(_13904_), .Y(_14656_) );
NAND2X1 NAND2X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_16598_), .B(_16600_), .Y(_14657_) );
XNOR2X1 XNOR2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_14657_), .B(bloque_datos[7]), .Y(_14658_) );
NOR2X1 NOR2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_14656_), .B(_14658_), .Y(_14659_) );
AND2X2 AND2X2_327 ( .gnd(gnd), .vdd(vdd), .A(_14658_), .B(_14656_), .Y(_14660_) );
NOR2X1 NOR2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_14659_), .B(_14660_), .Y(_14661_) );
NOR2X1 NOR2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_14651_), .B(_14661_), .Y(_14662_) );
AND2X2 AND2X2_328 ( .gnd(gnd), .vdd(vdd), .A(_14661_), .B(_14651_), .Y(_14663_) );
OAI21X1 OAI21X1_2306 ( .gnd(gnd), .vdd(vdd), .A(_14663_), .B(_14662_), .C(_14487_), .Y(_14664_) );
OR2X2 OR2X2_353 ( .gnd(gnd), .vdd(vdd), .A(_14661_), .B(_14651_), .Y(_14665_) );
NAND2X1 NAND2X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_14651_), .B(_14661_), .Y(_14666_) );
NAND3X1 NAND3X1_3305 ( .gnd(gnd), .vdd(vdd), .A(_14489_), .B(_14666_), .C(_14665_), .Y(_14667_) );
AND2X2 AND2X2_329 ( .gnd(gnd), .vdd(vdd), .A(_14667_), .B(_14664_), .Y(_14668_) );
AOI21X1 AOI21X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_13929_), .B(_13928_), .C(_13927_), .Y(_14669_) );
OAI21X1 OAI21X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_16617_), .B(_16612_), .C(bloque_datos_23_bF_buf3_), .Y(_14670_) );
NAND2X1 NAND2X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_16614_), .B(_16613_), .Y(_14671_) );
OR2X2 OR2X2_354 ( .gnd(gnd), .vdd(vdd), .A(_14671_), .B(bloque_datos_23_bF_buf2_), .Y(_14672_) );
NAND3X1 NAND3X1_3306 ( .gnd(gnd), .vdd(vdd), .A(_14670_), .B(_14669_), .C(_14672_), .Y(_14673_) );
INVX1 INVX1_2058 ( .gnd(gnd), .vdd(vdd), .A(_14670_), .Y(_14674_) );
NOR2X1 NOR2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf1_), .B(_14671_), .Y(_14675_) );
OAI21X1 OAI21X1_2308 ( .gnd(gnd), .vdd(vdd), .A(_14675_), .B(_14674_), .C(_13926_), .Y(_14676_) );
AOI21X1 AOI21X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_14673_), .B(_14676_), .C(_14668_), .Y(_14677_) );
NAND2X1 NAND2X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_14664_), .B(_14667_), .Y(_14678_) );
NAND2X1 NAND2X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_14676_), .B(_14673_), .Y(_14679_) );
NOR2X1 NOR2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_14678_), .B(_14679_), .Y(_14680_) );
OAI21X1 OAI21X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_14680_), .B(_14677_), .C(_14649_), .Y(_14681_) );
INVX1 INVX1_2059 ( .gnd(gnd), .vdd(vdd), .A(_14649_), .Y(_14682_) );
NOR3X1 NOR3X1_424 ( .gnd(gnd), .vdd(vdd), .A(_14675_), .B(_14674_), .C(_13926_), .Y(_14683_) );
AOI21X1 AOI21X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_14670_), .B(_14672_), .C(_14669_), .Y(_14684_) );
OAI21X1 OAI21X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_14683_), .B(_14684_), .C(_14678_), .Y(_14685_) );
NAND3X1 NAND3X1_3307 ( .gnd(gnd), .vdd(vdd), .A(_14673_), .B(_14676_), .C(_14668_), .Y(_14686_) );
NAND3X1 NAND3X1_3308 ( .gnd(gnd), .vdd(vdd), .A(_14685_), .B(_14686_), .C(_14682_), .Y(_14687_) );
NAND3X1 NAND3X1_3309 ( .gnd(gnd), .vdd(vdd), .A(_14495_), .B(_14687_), .C(_14681_), .Y(_14688_) );
OAI21X1 OAI21X1_2311 ( .gnd(gnd), .vdd(vdd), .A(_14680_), .B(_14677_), .C(_14682_), .Y(_14689_) );
NAND3X1 NAND3X1_3310 ( .gnd(gnd), .vdd(vdd), .A(_14649_), .B(_14685_), .C(_14686_), .Y(_14690_) );
NAND3X1 NAND3X1_3311 ( .gnd(gnd), .vdd(vdd), .A(_14500_), .B(_14690_), .C(_14689_), .Y(_14691_) );
NAND2X1 NAND2X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_14691_), .B(_14688_), .Y(_14692_) );
NAND2X1 NAND2X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_16631_), .B(_16630_), .Y(_14693_) );
XNOR2X1 XNOR2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_14693_), .B(bloque_datos[39]), .Y(_14694_) );
NOR2X1 NOR2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_13964_), .B(_14694_), .Y(_14695_) );
AND2X2 AND2X2_330 ( .gnd(gnd), .vdd(vdd), .A(_14694_), .B(_13964_), .Y(_14696_) );
OAI21X1 OAI21X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_14696_), .B(_14695_), .C(_14692_), .Y(_14697_) );
AND2X2 AND2X2_331 ( .gnd(gnd), .vdd(vdd), .A(_14688_), .B(_14691_), .Y(_14698_) );
OR2X2 OR2X2_355 ( .gnd(gnd), .vdd(vdd), .A(_14694_), .B(_13964_), .Y(_14699_) );
NAND2X1 NAND2X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_13964_), .B(_14694_), .Y(_14700_) );
NAND3X1 NAND3X1_3312 ( .gnd(gnd), .vdd(vdd), .A(_14699_), .B(_14700_), .C(_14698_), .Y(_14701_) );
NAND3X1 NAND3X1_3313 ( .gnd(gnd), .vdd(vdd), .A(_14648_), .B(_14697_), .C(_14701_), .Y(_14702_) );
OAI21X1 OAI21X1_2313 ( .gnd(gnd), .vdd(vdd), .A(_13974_), .B(_13976_), .C(_13969_), .Y(_14703_) );
AOI21X1 AOI21X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_14699_), .B(_14700_), .C(_14698_), .Y(_14704_) );
NOR3X1 NOR3X1_425 ( .gnd(gnd), .vdd(vdd), .A(_14695_), .B(_14696_), .C(_14692_), .Y(_14705_) );
OAI21X1 OAI21X1_2314 ( .gnd(gnd), .vdd(vdd), .A(_14704_), .B(_14705_), .C(_14703_), .Y(_14706_) );
NAND3X1 NAND3X1_3314 ( .gnd(gnd), .vdd(vdd), .A(_14510_), .B(_14702_), .C(_14706_), .Y(_14707_) );
NAND3X1 NAND3X1_3315 ( .gnd(gnd), .vdd(vdd), .A(_14703_), .B(_14697_), .C(_14701_), .Y(_14708_) );
OAI21X1 OAI21X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_14704_), .B(_14705_), .C(_14648_), .Y(_14709_) );
NAND3X1 NAND3X1_3316 ( .gnd(gnd), .vdd(vdd), .A(_14512_), .B(_14708_), .C(_14709_), .Y(_14710_) );
AND2X2 AND2X2_332 ( .gnd(gnd), .vdd(vdd), .A(_14707_), .B(_14710_), .Y(_14711_) );
XNOR2X1 XNOR2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_16640_), .B(bloque_datos[55]), .Y(_14712_) );
OR2X2 OR2X2_356 ( .gnd(gnd), .vdd(vdd), .A(_14712_), .B(_13999_), .Y(_14713_) );
NAND2X1 NAND2X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_13999_), .B(_14712_), .Y(_14714_) );
AOI21X1 AOI21X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_14714_), .B(_14713_), .C(_14711_), .Y(_14715_) );
NAND2X1 NAND2X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_14707_), .B(_14710_), .Y(_14716_) );
NOR2X1 NOR2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_13999_), .B(_14712_), .Y(_14717_) );
AND2X2 AND2X2_333 ( .gnd(gnd), .vdd(vdd), .A(_14712_), .B(_13999_), .Y(_14718_) );
NOR3X1 NOR3X1_426 ( .gnd(gnd), .vdd(vdd), .A(_14718_), .B(_14717_), .C(_14716_), .Y(_14719_) );
OAI21X1 OAI21X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_14715_), .B(_14719_), .C(_14647_), .Y(_14720_) );
OAI21X1 OAI21X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_14009_), .B(_14011_), .C(_14004_), .Y(_14721_) );
OAI21X1 OAI21X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_14718_), .B(_14717_), .C(_14716_), .Y(_14722_) );
NAND3X1 NAND3X1_3317 ( .gnd(gnd), .vdd(vdd), .A(_14714_), .B(_14713_), .C(_14711_), .Y(_14723_) );
NAND3X1 NAND3X1_3318 ( .gnd(gnd), .vdd(vdd), .A(_14722_), .B(_14721_), .C(_14723_), .Y(_14724_) );
NAND3X1 NAND3X1_3319 ( .gnd(gnd), .vdd(vdd), .A(_14646_), .B(_14724_), .C(_14720_), .Y(_14725_) );
OAI21X1 OAI21X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_14715_), .B(_14719_), .C(_14721_), .Y(_14726_) );
NAND3X1 NAND3X1_3320 ( .gnd(gnd), .vdd(vdd), .A(_14647_), .B(_14722_), .C(_14723_), .Y(_14727_) );
NAND3X1 NAND3X1_3321 ( .gnd(gnd), .vdd(vdd), .A(_14645_), .B(_14727_), .C(_14726_), .Y(_14728_) );
AND2X2 AND2X2_334 ( .gnd(gnd), .vdd(vdd), .A(_14725_), .B(_14728_), .Y(_14729_) );
OAI21X1 OAI21X1_2320 ( .gnd(gnd), .vdd(vdd), .A(_16646_), .B(_16652_), .C(bloque_datos_71_bF_buf3_), .Y(_14730_) );
INVX1 INVX1_2060 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf2_), .Y(_14731_) );
OAI21X1 OAI21X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_16648_), .B(_16651_), .C(_16647_), .Y(_14732_) );
NAND3X1 NAND3X1_3322 ( .gnd(gnd), .vdd(vdd), .A(_16577_), .B(_16645_), .C(_16642_), .Y(_14733_) );
NAND3X1 NAND3X1_3323 ( .gnd(gnd), .vdd(vdd), .A(_14731_), .B(_14732_), .C(_14733_), .Y(_14734_) );
NAND2X1 NAND2X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_14734_), .B(_14730_), .Y(_14735_) );
OR2X2 OR2X2_357 ( .gnd(gnd), .vdd(vdd), .A(_14735_), .B(_14037_), .Y(_14736_) );
NAND2X1 NAND2X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_14037_), .B(_14735_), .Y(_14737_) );
AOI21X1 AOI21X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_14736_), .B(_14737_), .C(_14729_), .Y(_14738_) );
NAND2X1 NAND2X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_14725_), .B(_14728_), .Y(_14739_) );
NOR2X1 NOR2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_14037_), .B(_14735_), .Y(_14740_) );
AND2X2 AND2X2_335 ( .gnd(gnd), .vdd(vdd), .A(_14735_), .B(_14037_), .Y(_14741_) );
NOR3X1 NOR3X1_427 ( .gnd(gnd), .vdd(vdd), .A(_14741_), .B(_14740_), .C(_14739_), .Y(_14742_) );
OAI21X1 OAI21X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_14738_), .B(_14742_), .C(_14644_), .Y(_14743_) );
AOI21X1 AOI21X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_14045_), .B(_13885_), .C(_14048_), .Y(_14744_) );
OAI21X1 OAI21X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_14741_), .B(_14740_), .C(_14739_), .Y(_14745_) );
NAND3X1 NAND3X1_3324 ( .gnd(gnd), .vdd(vdd), .A(_14736_), .B(_14737_), .C(_14729_), .Y(_14746_) );
NAND3X1 NAND3X1_3325 ( .gnd(gnd), .vdd(vdd), .A(_14744_), .B(_14745_), .C(_14746_), .Y(_14747_) );
AOI21X1 AOI21X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_14747_), .B(_14743_), .C(_14643_), .Y(_14748_) );
INVX1 INVX1_2061 ( .gnd(gnd), .vdd(vdd), .A(_14643_), .Y(_14749_) );
OAI21X1 OAI21X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_14738_), .B(_14742_), .C(_14744_), .Y(_14750_) );
NAND3X1 NAND3X1_3326 ( .gnd(gnd), .vdd(vdd), .A(_14745_), .B(_14644_), .C(_14746_), .Y(_14751_) );
AOI21X1 AOI21X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_14751_), .B(_14750_), .C(_14749_), .Y(_14752_) );
OR2X2 OR2X2_358 ( .gnd(gnd), .vdd(vdd), .A(_14748_), .B(_14752_), .Y(_14753_) );
NAND3X1 NAND3X1_3327 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf0_), .B(_16662_), .C(_16666_), .Y(_14754_) );
INVX1 INVX1_2062 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf3_), .Y(_14755_) );
OAI21X1 OAI21X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_16663_), .B(_16661_), .C(_14755_), .Y(_14756_) );
NAND2X1 NAND2X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_14754_), .B(_14756_), .Y(_14757_) );
OR2X2 OR2X2_359 ( .gnd(gnd), .vdd(vdd), .A(_14757_), .B(_14079_), .Y(_14758_) );
NAND2X1 NAND2X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_14079_), .B(_14757_), .Y(_14759_) );
NAND3X1 NAND3X1_3328 ( .gnd(gnd), .vdd(vdd), .A(_14758_), .B(_14759_), .C(_14753_), .Y(_14760_) );
NOR2X1 NOR2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_14748_), .B(_14752_), .Y(_14761_) );
NOR2X1 NOR2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_14079_), .B(_14757_), .Y(_14762_) );
AND2X2 AND2X2_336 ( .gnd(gnd), .vdd(vdd), .A(_14757_), .B(_14079_), .Y(_14763_) );
OAI21X1 OAI21X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_14763_), .B(_14762_), .C(_14761_), .Y(_14764_) );
NAND3X1 NAND3X1_3329 ( .gnd(gnd), .vdd(vdd), .A(_14764_), .B(_14642_), .C(_14760_), .Y(_14765_) );
AOI21X1 AOI21X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_14087_), .B(_13883_), .C(_14090_), .Y(_14766_) );
NOR3X1 NOR3X1_428 ( .gnd(gnd), .vdd(vdd), .A(_14763_), .B(_14762_), .C(_14761_), .Y(_14767_) );
AOI21X1 AOI21X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_14759_), .B(_14758_), .C(_14753_), .Y(_14768_) );
OAI21X1 OAI21X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_14767_), .B(_14768_), .C(_14766_), .Y(_14769_) );
AOI21X1 AOI21X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_14765_), .B(_14769_), .C(_14641_), .Y(_14770_) );
INVX1 INVX1_2063 ( .gnd(gnd), .vdd(vdd), .A(_14641_), .Y(_14771_) );
NAND3X1 NAND3X1_3330 ( .gnd(gnd), .vdd(vdd), .A(_14766_), .B(_14764_), .C(_14760_), .Y(_14772_) );
OAI21X1 OAI21X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_14767_), .B(_14768_), .C(_14642_), .Y(_14773_) );
AOI21X1 AOI21X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_14772_), .B(_14773_), .C(_14771_), .Y(_14774_) );
NOR2X1 NOR2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_14770_), .B(_14774_), .Y(_14775_) );
NAND3X1 NAND3X1_3331 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_135_), .B(_16674_), .C(_16677_), .Y(_14776_) );
INVX1 INVX1_2064 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_135_), .Y(_14777_) );
OAI21X1 OAI21X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_16675_), .B(_16673_), .C(_14777_), .Y(_14778_) );
NAND2X1 NAND2X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_14776_), .B(_14778_), .Y(_14779_) );
NOR2X1 NOR2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_14779_), .B(_14120_), .Y(_14780_) );
NAND2X1 NAND2X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_14779_), .B(_14120_), .Y(_14781_) );
INVX1 INVX1_2065 ( .gnd(gnd), .vdd(vdd), .A(_14781_), .Y(_14782_) );
NOR3X1 NOR3X1_429 ( .gnd(gnd), .vdd(vdd), .A(_14782_), .B(_14780_), .C(_14775_), .Y(_14783_) );
OR2X2 OR2X2_360 ( .gnd(gnd), .vdd(vdd), .A(_14770_), .B(_14774_), .Y(_14784_) );
INVX1 INVX1_2066 ( .gnd(gnd), .vdd(vdd), .A(_14780_), .Y(_14785_) );
AOI21X1 AOI21X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_14781_), .B(_14785_), .C(_14784_), .Y(_14786_) );
OAI21X1 OAI21X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_14783_), .B(_14786_), .C(_14640_), .Y(_14787_) );
NAND3X1 NAND3X1_3332 ( .gnd(gnd), .vdd(vdd), .A(_14781_), .B(_14785_), .C(_14784_), .Y(_14788_) );
OAI21X1 OAI21X1_2331 ( .gnd(gnd), .vdd(vdd), .A(_14782_), .B(_14780_), .C(_14775_), .Y(_14789_) );
NAND3X1 NAND3X1_3333 ( .gnd(gnd), .vdd(vdd), .A(_14639_), .B(_14789_), .C(_14788_), .Y(_14790_) );
AOI21X1 AOI21X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_14790_), .B(_14787_), .C(_14554_), .Y(_14791_) );
INVX1 INVX1_2067 ( .gnd(gnd), .vdd(vdd), .A(_14554_), .Y(_14792_) );
OAI21X1 OAI21X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_14783_), .B(_14786_), .C(_14639_), .Y(_14793_) );
NAND3X1 NAND3X1_3334 ( .gnd(gnd), .vdd(vdd), .A(_14789_), .B(_14788_), .C(_14640_), .Y(_14794_) );
AOI21X1 AOI21X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_14794_), .B(_14793_), .C(_14792_), .Y(_14795_) );
OAI21X1 OAI21X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_14791_), .B(_14795_), .C(_14638_), .Y(_14796_) );
NAND3X1 NAND3X1_3335 ( .gnd(gnd), .vdd(vdd), .A(_14792_), .B(_14794_), .C(_14793_), .Y(_14797_) );
NAND3X1 NAND3X1_3336 ( .gnd(gnd), .vdd(vdd), .A(_14554_), .B(_14790_), .C(_14787_), .Y(_14798_) );
NAND3X1 NAND3X1_3337 ( .gnd(gnd), .vdd(vdd), .A(_14160_), .B(_14797_), .C(_14798_), .Y(_14799_) );
NAND2X1 NAND2X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_14799_), .B(_14796_), .Y(_14800_) );
OAI21X1 OAI21X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_14171_), .B(_14193_), .C(_14800_), .Y(_14801_) );
INVX1 INVX1_2068 ( .gnd(gnd), .vdd(vdd), .A(_16686_), .Y(_14802_) );
OAI21X1 OAI21X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_14170_), .B(_14172_), .C(_14165_), .Y(_14803_) );
INVX1 INVX1_2069 ( .gnd(gnd), .vdd(vdd), .A(_14803_), .Y(_14804_) );
AND2X2 AND2X2_337 ( .gnd(gnd), .vdd(vdd), .A(_14796_), .B(_14799_), .Y(_14805_) );
AOI22X1 AOI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_16683_), .B(_14802_), .C(_14805_), .D(_14804_), .Y(_14806_) );
NAND3X1 NAND3X1_3338 ( .gnd(gnd), .vdd(vdd), .A(_14563_), .B(_14801_), .C(_14806_), .Y(_14807_) );
INVX1 INVX1_2070 ( .gnd(gnd), .vdd(vdd), .A(_14563_), .Y(_14808_) );
NOR2X1 NOR2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_14804_), .B(_14805_), .Y(_14809_) );
NAND2X1 NAND2X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_16683_), .B(_14802_), .Y(_14810_) );
OAI21X1 OAI21X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_14800_), .B(_14803_), .C(_14810_), .Y(_14811_) );
OAI21X1 OAI21X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_14809_), .B(_14811_), .C(_14808_), .Y(_14812_) );
AND2X2 AND2X2_338 ( .gnd(gnd), .vdd(vdd), .A(_14807_), .B(_14812_), .Y(_14813_) );
INVX1 INVX1_2071 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_151_), .Y(_14814_) );
AOI21X1 AOI21X1_2071 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_150_), .B(_14196_), .C(_14814_), .Y(_14815_) );
NOR3X1 NOR3X1_430 ( .gnd(gnd), .vdd(vdd), .A(_14198_), .B(module_3_W_151_), .C(_14201_), .Y(_14816_) );
OAI21X1 OAI21X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_14815_), .B(_14816_), .C(_14813_), .Y(_14817_) );
NAND2X1 NAND2X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_14812_), .B(_14807_), .Y(_14818_) );
OAI21X1 OAI21X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_14201_), .B(_14198_), .C(module_3_W_151_), .Y(_14819_) );
NAND3X1 NAND3X1_3339 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_150_), .B(_14814_), .C(_14196_), .Y(_14820_) );
NAND3X1 NAND3X1_3340 ( .gnd(gnd), .vdd(vdd), .A(_14819_), .B(_14820_), .C(_14818_), .Y(_14821_) );
AND2X2 AND2X2_339 ( .gnd(gnd), .vdd(vdd), .A(_14817_), .B(_14821_), .Y(_14822_) );
OAI21X1 OAI21X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_14227_), .B(_14207_), .C(_14822_), .Y(_14823_) );
OAI21X1 OAI21X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_13875_), .B(_14228_), .C(_14210_), .Y(_14824_) );
INVX1 INVX1_2072 ( .gnd(gnd), .vdd(vdd), .A(_14824_), .Y(_14825_) );
NAND2X1 NAND2X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_14821_), .B(_14817_), .Y(_14826_) );
AOI21X1 AOI21X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_14826_), .B(_14825_), .C(_16698_), .Y(_14827_) );
NAND3X1 NAND3X1_3341 ( .gnd(gnd), .vdd(vdd), .A(_14637_), .B(_14823_), .C(_14827_), .Y(_14828_) );
NOR2X1 NOR2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_14826_), .B(_14825_), .Y(_14829_) );
INVX1 INVX1_2073 ( .gnd(gnd), .vdd(vdd), .A(_16698_), .Y(_14830_) );
OAI21X1 OAI21X1_2342 ( .gnd(gnd), .vdd(vdd), .A(_14822_), .B(_14824_), .C(_14830_), .Y(_14831_) );
OAI21X1 OAI21X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_14831_), .B(_14829_), .C(_14576_), .Y(_14832_) );
NAND2X1 NAND2X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_14828_), .B(_14832_), .Y(_14833_) );
AOI21X1 AOI21X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_14634_), .B(_14636_), .C(_14833_), .Y(_14834_) );
NAND3X1 NAND3X1_3342 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_166_), .B(module_3_W_167_), .C(_14231_), .Y(_14835_) );
OAI21X1 OAI21X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_14236_), .B(_14233_), .C(_14635_), .Y(_14836_) );
AOI22X1 AOI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_14828_), .B(_14832_), .C(_14836_), .D(_14835_), .Y(_14837_) );
NOR2X1 NOR2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_14837_), .B(_14834_), .Y(_14838_) );
OAI21X1 OAI21X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_14262_), .B(_14242_), .C(_14838_), .Y(_14839_) );
OAI21X1 OAI21X1_2346 ( .gnd(gnd), .vdd(vdd), .A(_14263_), .B(_13873_), .C(_14245_), .Y(_14840_) );
INVX1 INVX1_2074 ( .gnd(gnd), .vdd(vdd), .A(_14840_), .Y(_14841_) );
NAND2X1 NAND2X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_14835_), .B(_14836_), .Y(_14842_) );
XNOR2X1 XNOR2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_14842_), .B(_14833_), .Y(_14843_) );
AOI22X1 AOI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_16706_), .B(_16708_), .C(_14843_), .D(_14841_), .Y(_14844_) );
NAND3X1 NAND3X1_3343 ( .gnd(gnd), .vdd(vdd), .A(_14633_), .B(_14839_), .C(_14844_), .Y(_14845_) );
NOR2X1 NOR2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_14843_), .B(_14841_), .Y(_14846_) );
OAI21X1 OAI21X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_14838_), .B(_14840_), .C(_16709_), .Y(_14847_) );
OAI21X1 OAI21X1_2348 ( .gnd(gnd), .vdd(vdd), .A(_14846_), .B(_14847_), .C(_14586_), .Y(_14848_) );
AND2X2 AND2X2_340 ( .gnd(gnd), .vdd(vdd), .A(_14845_), .B(_14848_), .Y(_14849_) );
INVX1 INVX1_2075 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_183_), .Y(_14850_) );
AOI21X1 AOI21X1_2074 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_182_), .B(_14266_), .C(_14850_), .Y(_14851_) );
NOR3X1 NOR3X1_431 ( .gnd(gnd), .vdd(vdd), .A(_14268_), .B(module_3_W_183_), .C(_14271_), .Y(_14852_) );
OAI21X1 OAI21X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_14851_), .B(_14852_), .C(_14849_), .Y(_14853_) );
NAND2X1 NAND2X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_14848_), .B(_14845_), .Y(_14854_) );
OAI21X1 OAI21X1_2350 ( .gnd(gnd), .vdd(vdd), .A(_14271_), .B(_14268_), .C(module_3_W_183_), .Y(_14855_) );
NAND3X1 NAND3X1_3344 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_182_), .B(_14850_), .C(_14266_), .Y(_14856_) );
NAND3X1 NAND3X1_3345 ( .gnd(gnd), .vdd(vdd), .A(_14855_), .B(_14856_), .C(_14854_), .Y(_14857_) );
NAND2X1 NAND2X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_14857_), .B(_14853_), .Y(_14858_) );
NOR2X1 NOR2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_14858_), .B(_14632_), .Y(_14859_) );
AND2X2 AND2X2_341 ( .gnd(gnd), .vdd(vdd), .A(_14853_), .B(_14857_), .Y(_14860_) );
OAI21X1 OAI21X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_14860_), .B(_14631_), .C(_13291_), .Y(_14861_) );
OAI21X1 OAI21X1_2352 ( .gnd(gnd), .vdd(vdd), .A(_14861_), .B(_14859_), .C(module_3_W_199_), .Y(_14862_) );
INVX1 INVX1_2076 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_199_), .Y(_14863_) );
OAI21X1 OAI21X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_14281_), .B(_14300_), .C(_14860_), .Y(_14865_) );
AOI21X1 AOI21X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_14858_), .B(_14632_), .C(_16723_), .Y(_14866_) );
NAND3X1 NAND3X1_3346 ( .gnd(gnd), .vdd(vdd), .A(_14863_), .B(_14865_), .C(_14866_), .Y(_14867_) );
NAND2X1 NAND2X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_14867_), .B(_14862_), .Y(_14868_) );
NOR3X1 NOR3X1_432 ( .gnd(gnd), .vdd(vdd), .A(_14300_), .B(_14302_), .C(_14301_), .Y(_14869_) );
NOR3X1 NOR3X1_433 ( .gnd(gnd), .vdd(vdd), .A(_13867_), .B(_14307_), .C(_14869_), .Y(_14870_) );
OAI21X1 OAI21X1_2354 ( .gnd(gnd), .vdd(vdd), .A(_14870_), .B(_14306_), .C(_14595_), .Y(_14871_) );
INVX2 INVX2_527 ( .gnd(gnd), .vdd(vdd), .A(_14595_), .Y(_14872_) );
NAND3X1 NAND3X1_3347 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_198_), .B(_14872_), .C(_14304_), .Y(_14873_) );
NAND3X1 NAND3X1_3348 ( .gnd(gnd), .vdd(vdd), .A(_14871_), .B(_14873_), .C(_14868_), .Y(_14874_) );
AND2X2 AND2X2_342 ( .gnd(gnd), .vdd(vdd), .A(_14862_), .B(_14867_), .Y(_14876_) );
AOI21X1 AOI21X1_2076 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_198_), .B(_14304_), .C(_14872_), .Y(_14877_) );
INVX1 INVX1_2077 ( .gnd(gnd), .vdd(vdd), .A(_14873_), .Y(_14878_) );
OAI21X1 OAI21X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_14878_), .B(_14877_), .C(_14876_), .Y(_14879_) );
AOI21X1 AOI21X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_14874_), .B(_14879_), .C(_14630_), .Y(_14880_) );
OAI21X1 OAI21X1_2356 ( .gnd(gnd), .vdd(vdd), .A(_14337_), .B(_13866_), .C(_14317_), .Y(_14881_) );
NAND2X1 NAND2X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_14874_), .B(_14879_), .Y(_14882_) );
OAI21X1 OAI21X1_2357 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .B(_14881_), .C(_16738_), .Y(_14883_) );
NOR3X1 NOR3X1_434 ( .gnd(gnd), .vdd(vdd), .A(_14880_), .B(_14606_), .C(_14883_), .Y(_14884_) );
INVX2 INVX2_528 ( .gnd(gnd), .vdd(vdd), .A(_14606_), .Y(_14885_) );
INVX1 INVX1_2078 ( .gnd(gnd), .vdd(vdd), .A(_14880_), .Y(_14887_) );
AND2X2 AND2X2_343 ( .gnd(gnd), .vdd(vdd), .A(_14879_), .B(_14874_), .Y(_14888_) );
AOI21X1 AOI21X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_14630_), .B(_14888_), .C(_16741_), .Y(_14889_) );
AOI21X1 AOI21X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_14887_), .B(_14889_), .C(_14885_), .Y(_14890_) );
NOR2X1 NOR2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_14884_), .B(_14890_), .Y(_14891_) );
INVX1 INVX1_2079 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_215_), .Y(_14892_) );
AOI21X1 AOI21X1_2080 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_214_), .B(_14340_), .C(_14892_), .Y(_14893_) );
NOR3X1 NOR3X1_435 ( .gnd(gnd), .vdd(vdd), .A(_14342_), .B(module_3_W_215_), .C(_14345_), .Y(_14894_) );
OAI21X1 OAI21X1_2358 ( .gnd(gnd), .vdd(vdd), .A(_14893_), .B(_14894_), .C(_14891_), .Y(_14895_) );
NAND3X1 NAND3X1_3349 ( .gnd(gnd), .vdd(vdd), .A(_14885_), .B(_14887_), .C(_14889_), .Y(_14896_) );
OAI21X1 OAI21X1_2359 ( .gnd(gnd), .vdd(vdd), .A(_14883_), .B(_14880_), .C(_14606_), .Y(_14898_) );
NAND2X1 NAND2X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_14898_), .B(_14896_), .Y(_14899_) );
OAI21X1 OAI21X1_2360 ( .gnd(gnd), .vdd(vdd), .A(_14345_), .B(_14342_), .C(module_3_W_215_), .Y(_14900_) );
NAND3X1 NAND3X1_3350 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_214_), .B(_14892_), .C(_14340_), .Y(_14901_) );
NAND3X1 NAND3X1_3351 ( .gnd(gnd), .vdd(vdd), .A(_14900_), .B(_14901_), .C(_14899_), .Y(_14902_) );
AND2X2 AND2X2_344 ( .gnd(gnd), .vdd(vdd), .A(_14895_), .B(_14902_), .Y(_14903_) );
OAI21X1 OAI21X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_14373_), .B(_14351_), .C(_14903_), .Y(_14904_) );
AOI21X1 AOI21X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_14355_), .B(_14353_), .C(_14373_), .Y(_14905_) );
NAND2X1 NAND2X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .B(_14895_), .Y(_14906_) );
AOI21X1 AOI21X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_14905_), .B(_14906_), .C(_16750_), .Y(_14907_) );
NAND3X1 NAND3X1_3352 ( .gnd(gnd), .vdd(vdd), .A(_14629_), .B(_14907_), .C(_14904_), .Y(_14909_) );
NOR2X1 NOR2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_14905_), .B(_14906_), .Y(_14910_) );
INVX1 INVX1_2080 ( .gnd(gnd), .vdd(vdd), .A(_16750_), .Y(_14911_) );
OAI21X1 OAI21X1_2362 ( .gnd(gnd), .vdd(vdd), .A(_14374_), .B(_13863_), .C(_14354_), .Y(_14912_) );
OAI21X1 OAI21X1_2363 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .B(_14912_), .C(_14911_), .Y(_14913_) );
OAI21X1 OAI21X1_2364 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .B(_14910_), .C(_14616_), .Y(_14914_) );
AND2X2 AND2X2_345 ( .gnd(gnd), .vdd(vdd), .A(_14914_), .B(_14909_), .Y(_14915_) );
INVX1 INVX1_2081 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_231_), .Y(_14916_) );
AOI21X1 AOI21X1_2083 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_230_), .B(_14377_), .C(_14916_), .Y(_14917_) );
NOR3X1 NOR3X1_436 ( .gnd(gnd), .vdd(vdd), .A(_14379_), .B(module_3_W_231_), .C(_14382_), .Y(_14918_) );
OAI21X1 OAI21X1_2365 ( .gnd(gnd), .vdd(vdd), .A(_14917_), .B(_14918_), .C(_14915_), .Y(_14920_) );
NAND2X1 NAND2X1_1958 ( .gnd(gnd), .vdd(vdd), .A(_14909_), .B(_14914_), .Y(_14921_) );
OAI21X1 OAI21X1_2366 ( .gnd(gnd), .vdd(vdd), .A(_14382_), .B(_14379_), .C(module_3_W_231_), .Y(_14922_) );
NAND3X1 NAND3X1_3353 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_230_), .B(_14916_), .C(_14377_), .Y(_14923_) );
NAND3X1 NAND3X1_3354 ( .gnd(gnd), .vdd(vdd), .A(_14922_), .B(_14923_), .C(_14921_), .Y(_14924_) );
AND2X2 AND2X2_346 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .B(_14924_), .Y(_14925_) );
OAI21X1 OAI21X1_2367 ( .gnd(gnd), .vdd(vdd), .A(_14410_), .B(_14388_), .C(_14925_), .Y(_14926_) );
OAI21X1 OAI21X1_2368 ( .gnd(gnd), .vdd(vdd), .A(_14411_), .B(_13857_), .C(_14391_), .Y(_14927_) );
INVX1 INVX1_2082 ( .gnd(gnd), .vdd(vdd), .A(_14927_), .Y(_14928_) );
NAND2X1 NAND2X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .B(_14920_), .Y(_14929_) );
AOI21X1 AOI21X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_14929_), .B(_14928_), .C(_16763_), .Y(_14931_) );
NAND3X1 NAND3X1_3355 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_247_), .B(_14926_), .C(_14931_), .Y(_14932_) );
INVX2 INVX2_529 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_247_), .Y(_14933_) );
NOR2X1 NOR2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_14929_), .B(_14928_), .Y(_14934_) );
INVX1 INVX1_2083 ( .gnd(gnd), .vdd(vdd), .A(_16763_), .Y(_14935_) );
OAI21X1 OAI21X1_2369 ( .gnd(gnd), .vdd(vdd), .A(_14925_), .B(_14927_), .C(_14935_), .Y(_14936_) );
OAI21X1 OAI21X1_2370 ( .gnd(gnd), .vdd(vdd), .A(_14936_), .B(_14934_), .C(_14933_), .Y(_14937_) );
NAND3X1 NAND3X1_3356 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .B(_14937_), .C(_14415_), .Y(_14938_) );
NOR2X1 NOR2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_14416_), .B(_14419_), .Y(_14939_) );
NOR3X1 NOR3X1_437 ( .gnd(gnd), .vdd(vdd), .A(_14934_), .B(_14933_), .C(_14936_), .Y(_14940_) );
AOI21X1 AOI21X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_14926_), .B(_14931_), .C(module_3_W_247_), .Y(_14942_) );
OAI21X1 OAI21X1_2371 ( .gnd(gnd), .vdd(vdd), .A(_14940_), .B(_14942_), .C(_14939_), .Y(_14943_) );
NAND3X1 NAND3X1_3357 ( .gnd(gnd), .vdd(vdd), .A(_14628_), .B(_14938_), .C(_14943_), .Y(_14944_) );
NAND3X1 NAND3X1_3358 ( .gnd(gnd), .vdd(vdd), .A(_14933_), .B(_14926_), .C(_14931_), .Y(_14945_) );
OAI21X1 OAI21X1_2372 ( .gnd(gnd), .vdd(vdd), .A(_14936_), .B(_14934_), .C(module_3_W_247_), .Y(_14946_) );
AOI22X1 AOI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_246_), .B(_14414_), .C(_14946_), .D(_14945_), .Y(_14947_) );
AOI21X1 AOI21X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .B(_14937_), .C(_14415_), .Y(_14948_) );
OAI21X1 OAI21X1_2373 ( .gnd(gnd), .vdd(vdd), .A(_14948_), .B(_14947_), .C(_14627_), .Y(_14949_) );
NAND3X1 NAND3X1_3359 ( .gnd(gnd), .vdd(vdd), .A(_14944_), .B(_14949_), .C(_14452_), .Y(_14950_) );
AOI21X1 AOI21X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_14415_), .B(_14420_), .C(_13832_), .Y(_14951_) );
OAI21X1 OAI21X1_2374 ( .gnd(gnd), .vdd(vdd), .A(_14951_), .B(_13855_), .C(_14427_), .Y(_14953_) );
NOR3X1 NOR3X1_438 ( .gnd(gnd), .vdd(vdd), .A(_14947_), .B(_14627_), .C(_14948_), .Y(_14954_) );
AOI21X1 AOI21X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_14938_), .B(_14943_), .C(_14628_), .Y(_14955_) );
OAI21X1 OAI21X1_2375 ( .gnd(gnd), .vdd(vdd), .A(_14954_), .B(_14955_), .C(_14953_), .Y(_14956_) );
NAND2X1 NAND2X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_14956_), .B(_14950_), .Y(_14957_) );
NAND2X1 NAND2X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_14957_), .B(_14450_), .Y(_14958_) );
OAI21X1 OAI21X1_2376 ( .gnd(gnd), .vdd(vdd), .A(_14954_), .B(_14955_), .C(_14452_), .Y(_14959_) );
NAND3X1 NAND3X1_3360 ( .gnd(gnd), .vdd(vdd), .A(_14944_), .B(_14949_), .C(_14953_), .Y(_14960_) );
NAND2X1 NAND2X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_14960_), .B(_14959_), .Y(_14961_) );
NAND3X1 NAND3X1_3361 ( .gnd(gnd), .vdd(vdd), .A(_13854_), .B(_14961_), .C(_14447_), .Y(_14962_) );
NAND2X1 NAND2X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_14962_), .B(_14958_), .Y(module_3_H_7_) );
NOR2X1 NOR2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_248_), .B(_13379_), .Y(_14964_) );
INVX1 INVX1_2084 ( .gnd(gnd), .vdd(vdd), .A(_14964_), .Y(_14965_) );
OAI21X1 OAI21X1_2377 ( .gnd(gnd), .vdd(vdd), .A(_13374_), .B(_13373_), .C(module_3_W_248_), .Y(_14966_) );
NAND2X1 NAND2X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_14966_), .B(_14965_), .Y(module_3_H_16_) );
XNOR2X1 XNOR2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_13506_), .B(module_3_W_249_), .Y(_14967_) );
INVX1 INVX1_2085 ( .gnd(gnd), .vdd(vdd), .A(_14967_), .Y(_14968_) );
OAI21X1 OAI21X1_2378 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_248_), .B(_13379_), .C(_14968_), .Y(_14969_) );
INVX2 INVX2_530 ( .gnd(gnd), .vdd(vdd), .A(_14969_), .Y(_14970_) );
NOR2X1 NOR2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_14965_), .B(_14968_), .Y(_14971_) );
NOR2X1 NOR2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_14971_), .B(_14970_), .Y(module_3_H_17_) );
NOR2X1 NOR2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_249_), .B(_13849_), .Y(_14973_) );
INVX1 INVX1_2086 ( .gnd(gnd), .vdd(vdd), .A(_14973_), .Y(_14974_) );
NAND2X1 NAND2X1_1965 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_250_), .B(_14441_), .Y(_14975_) );
OR2X2 OR2X2_361 ( .gnd(gnd), .vdd(vdd), .A(_14441_), .B(module_3_W_250_), .Y(_14976_) );
AOI21X1 AOI21X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_14975_), .B(_14976_), .C(_14974_), .Y(_14977_) );
INVX1 INVX1_2087 ( .gnd(gnd), .vdd(vdd), .A(_14977_), .Y(_14978_) );
NAND3X1 NAND3X1_3362 ( .gnd(gnd), .vdd(vdd), .A(_14974_), .B(_14975_), .C(_14976_), .Y(_14979_) );
NAND2X1 NAND2X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_14979_), .B(_14978_), .Y(_14980_) );
XNOR2X1 XNOR2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_14980_), .B(_14970_), .Y(module_3_H_18_) );
OAI21X1 OAI21X1_2379 ( .gnd(gnd), .vdd(vdd), .A(_14977_), .B(_14969_), .C(_14979_), .Y(_14982_) );
NOR2X1 NOR2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_250_), .B(_14442_), .Y(_14983_) );
INVX1 INVX1_2088 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_251_), .Y(_14984_) );
OAI21X1 OAI21X1_2380 ( .gnd(gnd), .vdd(vdd), .A(_14626_), .B(_14623_), .C(_14984_), .Y(_14985_) );
NAND2X1 NAND2X1_1967 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_251_), .B(_14627_), .Y(_14986_) );
NAND3X1 NAND3X1_3363 ( .gnd(gnd), .vdd(vdd), .A(_14983_), .B(_14985_), .C(_14986_), .Y(_14987_) );
AOI21X1 AOI21X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_14985_), .B(_14986_), .C(_14983_), .Y(_14988_) );
INVX1 INVX1_2089 ( .gnd(gnd), .vdd(vdd), .A(_14988_), .Y(_14989_) );
NAND2X1 NAND2X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_14987_), .B(_14989_), .Y(_14990_) );
XNOR2X1 XNOR2X1_389 ( .gnd(gnd), .vdd(vdd), .A(_14990_), .B(_14982_), .Y(module_3_H_19_) );
AOI21X1 AOI21X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_14982_), .B(_14987_), .C(_14988_), .Y(_14992_) );
OAI21X1 OAI21X1_2381 ( .gnd(gnd), .vdd(vdd), .A(_14453_), .B(_14621_), .C(_14619_), .Y(_14993_) );
INVX2 INVX2_531 ( .gnd(gnd), .vdd(vdd), .A(_14618_), .Y(_14994_) );
OAI21X1 OAI21X1_2382 ( .gnd(gnd), .vdd(vdd), .A(_14608_), .B(_14607_), .C(_14398_), .Y(_14995_) );
AOI21X1 AOI21X1_2092 ( .gnd(gnd), .vdd(vdd), .A(_14995_), .B(_14454_), .C(_14609_), .Y(_14996_) );
NOR3X1 NOR3X1_439 ( .gnd(gnd), .vdd(vdd), .A(_14361_), .B(_14597_), .C(_14600_), .Y(_14997_) );
AOI21X1 AOI21X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_14601_), .B(_14604_), .C(_14997_), .Y(_14998_) );
OAI21X1 OAI21X1_2383 ( .gnd(gnd), .vdd(vdd), .A(_14593_), .B(_14590_), .C(_14588_), .Y(_14999_) );
INVX1 INVX1_2090 ( .gnd(gnd), .vdd(vdd), .A(_14587_), .Y(_15000_) );
OR2X2 OR2X2_362 ( .gnd(gnd), .vdd(vdd), .A(_14578_), .B(_14461_), .Y(_15001_) );
OAI21X1 OAI21X1_2384 ( .gnd(gnd), .vdd(vdd), .A(_14580_), .B(_14459_), .C(_15001_), .Y(_15003_) );
NOR2X1 NOR2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_14462_), .B(_14637_), .Y(_15004_) );
OAI21X1 OAI21X1_2385 ( .gnd(gnd), .vdd(vdd), .A(_14565_), .B(_14566_), .C(_14251_), .Y(_15005_) );
AOI21X1 AOI21X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_15005_), .B(_14463_), .C(_14567_), .Y(_15006_) );
OAI21X1 OAI21X1_2386 ( .gnd(gnd), .vdd(vdd), .A(_14561_), .B(_14465_), .C(_14557_), .Y(_15007_) );
INVX2 INVX2_532 ( .gnd(gnd), .vdd(vdd), .A(_15007_), .Y(_15008_) );
NAND2X1 NAND2X1_1969 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_139_), .B(_14554_), .Y(_15009_) );
AND2X2 AND2X2_347 ( .gnd(gnd), .vdd(vdd), .A(_14551_), .B(_14547_), .Y(_15010_) );
INVX1 INVX1_2091 ( .gnd(gnd), .vdd(vdd), .A(_14548_), .Y(_15011_) );
INVX1 INVX1_2092 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf3_), .Y(_15012_) );
XNOR2X1 XNOR2X1_390 ( .gnd(gnd), .vdd(vdd), .A(_13183_), .B(_15507_), .Y(_15014_) );
NAND2X1 NAND2X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_14536_), .B(_14541_), .Y(_15015_) );
XOR2X1 XOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_13158_), .B(_15035_), .Y(_15016_) );
INVX1 INVX1_2093 ( .gnd(gnd), .vdd(vdd), .A(_14470_), .Y(_15017_) );
AOI21X1 AOI21X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_14524_), .B(_14522_), .C(_14098_), .Y(_15018_) );
OAI21X1 OAI21X1_2387 ( .gnd(gnd), .vdd(vdd), .A(_15017_), .B(_15018_), .C(_14525_), .Y(_15019_) );
XNOR2X1 XNOR2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_13132_), .B(_15002_), .Y(_15020_) );
OAI21X1 OAI21X1_2388 ( .gnd(gnd), .vdd(vdd), .A(_14061_), .B(_13428_), .C(_14064_), .Y(_15021_) );
AOI21X1 AOI21X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_14515_), .B(_15021_), .C(_14514_), .Y(_15022_) );
INVX1 INVX1_2094 ( .gnd(gnd), .vdd(vdd), .A(_14511_), .Y(_15023_) );
INVX1 INVX1_2095 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf1_), .Y(_15025_) );
AOI21X1 AOI21X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_14508_), .B(_14506_), .C(_14503_), .Y(_15026_) );
NOR2X1 NOR2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf1_), .B(_14500_), .Y(_15027_) );
INVX1 INVX1_2096 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf3_), .Y(_15028_) );
XNOR2X1 XNOR2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_16893_), .B(_14941_), .Y(_15029_) );
INVX1 INVX1_2097 ( .gnd(gnd), .vdd(vdd), .A(_15029_), .Y(_15030_) );
OAI21X1 OAI21X1_2389 ( .gnd(gnd), .vdd(vdd), .A(_14494_), .B(_14476_), .C(_14492_), .Y(_15031_) );
XNOR2X1 XNOR2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_16869_), .B(_14919_), .Y(_15032_) );
INVX1 INVX1_2098 ( .gnd(gnd), .vdd(vdd), .A(_15032_), .Y(_15033_) );
AOI21X1 AOI21X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_13948_), .B(_13406_), .C(_13952_), .Y(_15034_) );
OAI21X1 OAI21X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_15034_), .B(_14486_), .C(_14484_), .Y(_15036_) );
INVX1 INVX1_2099 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_28_), .Y(_15037_) );
XNOR2X1 XNOR2X1_394 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_0_), .B(module_3_W_12_), .Y(_15038_) );
XOR2X1 XOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_15038_), .B(module_3_W_8_), .Y(_15039_) );
NAND2X1 NAND2X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_15037_), .B(_15039_), .Y(_15040_) );
XNOR2X1 XNOR2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_15038_), .B(module_3_W_8_), .Y(_15041_) );
NAND2X1 NAND2X1_1972 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_28_), .B(_15041_), .Y(_15042_) );
NAND3X1 NAND3X1_3364 ( .gnd(gnd), .vdd(vdd), .A(_14480_), .B(_15042_), .C(_15040_), .Y(_15043_) );
AOI21X1 AOI21X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_15042_), .B(_15040_), .C(_14480_), .Y(_15044_) );
INVX2 INVX2_533 ( .gnd(gnd), .vdd(vdd), .A(_15044_), .Y(_15045_) );
AOI21X1 AOI21X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_15043_), .B(_15045_), .C(_15036_), .Y(_15047_) );
INVX1 INVX1_2100 ( .gnd(gnd), .vdd(vdd), .A(_14484_), .Y(_15048_) );
AOI21X1 AOI21X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_14485_), .B(_14479_), .C(_15048_), .Y(_15049_) );
INVX2 INVX2_534 ( .gnd(gnd), .vdd(vdd), .A(_15043_), .Y(_15050_) );
NOR3X1 NOR3X1_440 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .B(_15044_), .C(_15050_), .Y(_15051_) );
OAI21X1 OAI21X1_2391 ( .gnd(gnd), .vdd(vdd), .A(_15051_), .B(_15047_), .C(_15033_), .Y(_15052_) );
OAI21X1 OAI21X1_2392 ( .gnd(gnd), .vdd(vdd), .A(_15050_), .B(_15044_), .C(_15049_), .Y(_15053_) );
NAND3X1 NAND3X1_3365 ( .gnd(gnd), .vdd(vdd), .A(_15036_), .B(_15043_), .C(_15045_), .Y(_15054_) );
NAND3X1 NAND3X1_3366 ( .gnd(gnd), .vdd(vdd), .A(_15032_), .B(_15054_), .C(_15053_), .Y(_15055_) );
NAND3X1 NAND3X1_3367 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf0_), .B(_15055_), .C(_15052_), .Y(_15056_) );
INVX1 INVX1_2101 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf3_), .Y(_15058_) );
NAND3X1 NAND3X1_3368 ( .gnd(gnd), .vdd(vdd), .A(_15033_), .B(_15054_), .C(_15053_), .Y(_15059_) );
OAI21X1 OAI21X1_2393 ( .gnd(gnd), .vdd(vdd), .A(_15051_), .B(_15047_), .C(_15032_), .Y(_15060_) );
NAND3X1 NAND3X1_3369 ( .gnd(gnd), .vdd(vdd), .A(_15058_), .B(_15059_), .C(_15060_), .Y(_15061_) );
NAND3X1 NAND3X1_3370 ( .gnd(gnd), .vdd(vdd), .A(_14488_), .B(_15056_), .C(_15061_), .Y(_15062_) );
INVX1 INVX1_2102 ( .gnd(gnd), .vdd(vdd), .A(_14488_), .Y(_15063_) );
NAND3X1 NAND3X1_3371 ( .gnd(gnd), .vdd(vdd), .A(_15058_), .B(_15055_), .C(_15052_), .Y(_15064_) );
NAND3X1 NAND3X1_3372 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf2_), .B(_15059_), .C(_15060_), .Y(_15065_) );
NAND3X1 NAND3X1_3373 ( .gnd(gnd), .vdd(vdd), .A(_15063_), .B(_15064_), .C(_15065_), .Y(_15066_) );
AOI21X1 AOI21X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .B(_15066_), .C(_15031_), .Y(_15067_) );
INVX1 INVX1_2103 ( .gnd(gnd), .vdd(vdd), .A(_14492_), .Y(_15069_) );
AOI21X1 AOI21X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_14493_), .B(_14499_), .C(_15069_), .Y(_15070_) );
AOI21X1 AOI21X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_15064_), .B(_15065_), .C(_15063_), .Y(_15071_) );
AOI21X1 AOI21X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_15056_), .B(_15061_), .C(_14488_), .Y(_15072_) );
NOR3X1 NOR3X1_441 ( .gnd(gnd), .vdd(vdd), .A(_15071_), .B(_15070_), .C(_15072_), .Y(_15073_) );
OAI21X1 OAI21X1_2394 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_15067_), .C(_15030_), .Y(_15074_) );
OAI21X1 OAI21X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_15071_), .B(_15072_), .C(_15070_), .Y(_15075_) );
NAND3X1 NAND3X1_3374 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .B(_15066_), .C(_15031_), .Y(_15076_) );
NAND3X1 NAND3X1_3375 ( .gnd(gnd), .vdd(vdd), .A(_15029_), .B(_15075_), .C(_15076_), .Y(_15077_) );
NAND3X1 NAND3X1_3376 ( .gnd(gnd), .vdd(vdd), .A(_15028_), .B(_15077_), .C(_15074_), .Y(_15078_) );
NAND3X1 NAND3X1_3377 ( .gnd(gnd), .vdd(vdd), .A(_15030_), .B(_15075_), .C(_15076_), .Y(_15080_) );
OAI21X1 OAI21X1_2396 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_15067_), .C(_15029_), .Y(_15081_) );
NAND3X1 NAND3X1_3378 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf2_), .B(_15080_), .C(_15081_), .Y(_15082_) );
AOI21X1 AOI21X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_15078_), .B(_15082_), .C(_15027_), .Y(_15083_) );
INVX1 INVX1_2104 ( .gnd(gnd), .vdd(vdd), .A(_15027_), .Y(_15084_) );
NAND3X1 NAND3X1_3379 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf1_), .B(_15077_), .C(_15074_), .Y(_15085_) );
NAND3X1 NAND3X1_3380 ( .gnd(gnd), .vdd(vdd), .A(_15028_), .B(_15080_), .C(_15081_), .Y(_15086_) );
AOI21X1 AOI21X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_15085_), .B(_15086_), .C(_15084_), .Y(_15087_) );
OAI21X1 OAI21X1_2397 ( .gnd(gnd), .vdd(vdd), .A(_15083_), .B(_15087_), .C(_15026_), .Y(_15088_) );
OAI21X1 OAI21X1_2398 ( .gnd(gnd), .vdd(vdd), .A(_14474_), .B(_14504_), .C(_14507_), .Y(_15089_) );
NAND3X1 NAND3X1_3381 ( .gnd(gnd), .vdd(vdd), .A(_15084_), .B(_15085_), .C(_15086_), .Y(_15091_) );
NAND3X1 NAND3X1_3382 ( .gnd(gnd), .vdd(vdd), .A(_15027_), .B(_15078_), .C(_15082_), .Y(_15092_) );
NAND3X1 NAND3X1_3383 ( .gnd(gnd), .vdd(vdd), .A(_15091_), .B(_15092_), .C(_15089_), .Y(_15093_) );
XNOR2X1 XNOR2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_13107_), .B(_14972_), .Y(_15094_) );
NAND3X1 NAND3X1_3384 ( .gnd(gnd), .vdd(vdd), .A(_15094_), .B(_15093_), .C(_15088_), .Y(_15095_) );
AOI21X1 AOI21X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_15091_), .B(_15092_), .C(_15089_), .Y(_15096_) );
NOR3X1 NOR3X1_442 ( .gnd(gnd), .vdd(vdd), .A(_15083_), .B(_15087_), .C(_15026_), .Y(_15097_) );
INVX1 INVX1_2105 ( .gnd(gnd), .vdd(vdd), .A(_15094_), .Y(_15098_) );
OAI21X1 OAI21X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_15097_), .B(_15096_), .C(_15098_), .Y(_15099_) );
NAND3X1 NAND3X1_3385 ( .gnd(gnd), .vdd(vdd), .A(_15025_), .B(_15095_), .C(_15099_), .Y(_15100_) );
NAND3X1 NAND3X1_3386 ( .gnd(gnd), .vdd(vdd), .A(_15098_), .B(_15093_), .C(_15088_), .Y(_15102_) );
OAI21X1 OAI21X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_15097_), .B(_15096_), .C(_15094_), .Y(_15103_) );
NAND3X1 NAND3X1_3387 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf0_), .B(_15102_), .C(_15103_), .Y(_15104_) );
AOI21X1 AOI21X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_15100_), .B(_15104_), .C(_15023_), .Y(_15105_) );
NAND3X1 NAND3X1_3388 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf4_), .B(_15095_), .C(_15099_), .Y(_15106_) );
NAND3X1 NAND3X1_3389 ( .gnd(gnd), .vdd(vdd), .A(_15025_), .B(_15102_), .C(_15103_), .Y(_15107_) );
AOI21X1 AOI21X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_15106_), .B(_15107_), .C(_14511_), .Y(_15108_) );
OAI21X1 OAI21X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_15105_), .B(_15108_), .C(_15022_), .Y(_15109_) );
INVX1 INVX1_2106 ( .gnd(gnd), .vdd(vdd), .A(_14514_), .Y(_15110_) );
OAI21X1 OAI21X1_2402 ( .gnd(gnd), .vdd(vdd), .A(_14471_), .B(_14516_), .C(_15110_), .Y(_15111_) );
NAND3X1 NAND3X1_3390 ( .gnd(gnd), .vdd(vdd), .A(_14511_), .B(_15106_), .C(_15107_), .Y(_15113_) );
NAND3X1 NAND3X1_3391 ( .gnd(gnd), .vdd(vdd), .A(_15023_), .B(_15100_), .C(_15104_), .Y(_15114_) );
NAND3X1 NAND3X1_3392 ( .gnd(gnd), .vdd(vdd), .A(_15113_), .B(_15114_), .C(_15111_), .Y(_15115_) );
NAND3X1 NAND3X1_3393 ( .gnd(gnd), .vdd(vdd), .A(_15020_), .B(_15109_), .C(_15115_), .Y(_15116_) );
INVX1 INVX1_2107 ( .gnd(gnd), .vdd(vdd), .A(_15020_), .Y(_15117_) );
AOI21X1 AOI21X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_15113_), .B(_15114_), .C(_15111_), .Y(_15118_) );
NOR3X1 NOR3X1_443 ( .gnd(gnd), .vdd(vdd), .A(_15105_), .B(_15108_), .C(_15022_), .Y(_15119_) );
OAI21X1 OAI21X1_2403 ( .gnd(gnd), .vdd(vdd), .A(_15119_), .B(_15118_), .C(_15117_), .Y(_15120_) );
NAND3X1 NAND3X1_3394 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf0_), .B(_15116_), .C(_15120_), .Y(_15121_) );
INVX1 INVX1_2108 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf3_), .Y(_15122_) );
NAND3X1 NAND3X1_3395 ( .gnd(gnd), .vdd(vdd), .A(_15117_), .B(_15109_), .C(_15115_), .Y(_15124_) );
OAI21X1 OAI21X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_15119_), .B(_15118_), .C(_15020_), .Y(_15125_) );
NAND3X1 NAND3X1_3396 ( .gnd(gnd), .vdd(vdd), .A(_15122_), .B(_15124_), .C(_15125_), .Y(_15126_) );
NAND3X1 NAND3X1_3397 ( .gnd(gnd), .vdd(vdd), .A(_14526_), .B(_15121_), .C(_15126_), .Y(_15127_) );
INVX1 INVX1_2109 ( .gnd(gnd), .vdd(vdd), .A(_14526_), .Y(_15128_) );
NAND3X1 NAND3X1_3398 ( .gnd(gnd), .vdd(vdd), .A(_15122_), .B(_15116_), .C(_15120_), .Y(_15129_) );
NAND3X1 NAND3X1_3399 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf2_), .B(_15124_), .C(_15125_), .Y(_15130_) );
NAND3X1 NAND3X1_3400 ( .gnd(gnd), .vdd(vdd), .A(_15128_), .B(_15129_), .C(_15130_), .Y(_15131_) );
AOI21X1 AOI21X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_15127_), .B(_15131_), .C(_15019_), .Y(_15132_) );
AOI21X1 AOI21X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_14527_), .B(_14526_), .C(_14101_), .Y(_15133_) );
AOI21X1 AOI21X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_14470_), .B(_14528_), .C(_15133_), .Y(_15135_) );
AOI21X1 AOI21X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_15129_), .B(_15130_), .C(_15128_), .Y(_15136_) );
AOI21X1 AOI21X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_15121_), .B(_15126_), .C(_14526_), .Y(_15137_) );
NOR3X1 NOR3X1_444 ( .gnd(gnd), .vdd(vdd), .A(_15136_), .B(_15137_), .C(_15135_), .Y(_15138_) );
OAI21X1 OAI21X1_2405 ( .gnd(gnd), .vdd(vdd), .A(_15138_), .B(_15132_), .C(_15016_), .Y(_15139_) );
INVX1 INVX1_2110 ( .gnd(gnd), .vdd(vdd), .A(_15016_), .Y(_15140_) );
OAI21X1 OAI21X1_2406 ( .gnd(gnd), .vdd(vdd), .A(_15136_), .B(_15137_), .C(_15135_), .Y(_15141_) );
NAND3X1 NAND3X1_3401 ( .gnd(gnd), .vdd(vdd), .A(_15127_), .B(_15131_), .C(_15019_), .Y(_15142_) );
NAND3X1 NAND3X1_3402 ( .gnd(gnd), .vdd(vdd), .A(_15140_), .B(_15141_), .C(_15142_), .Y(_15143_) );
NAND3X1 NAND3X1_3403 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf1_), .B(_15143_), .C(_15139_), .Y(_15144_) );
INVX1 INVX1_2111 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf0_), .Y(_15146_) );
NAND3X1 NAND3X1_3404 ( .gnd(gnd), .vdd(vdd), .A(_15016_), .B(_15141_), .C(_15142_), .Y(_15147_) );
OAI21X1 OAI21X1_2407 ( .gnd(gnd), .vdd(vdd), .A(_15138_), .B(_15132_), .C(_15140_), .Y(_15148_) );
NAND3X1 NAND3X1_3405 ( .gnd(gnd), .vdd(vdd), .A(_15146_), .B(_15147_), .C(_15148_), .Y(_15149_) );
NAND3X1 NAND3X1_3406 ( .gnd(gnd), .vdd(vdd), .A(_14537_), .B(_15144_), .C(_15149_), .Y(_15150_) );
INVX1 INVX1_2112 ( .gnd(gnd), .vdd(vdd), .A(_14537_), .Y(_15151_) );
NAND3X1 NAND3X1_3407 ( .gnd(gnd), .vdd(vdd), .A(_15146_), .B(_15143_), .C(_15139_), .Y(_15152_) );
NAND3X1 NAND3X1_3408 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf4_), .B(_15147_), .C(_15148_), .Y(_15153_) );
NAND3X1 NAND3X1_3409 ( .gnd(gnd), .vdd(vdd), .A(_15151_), .B(_15152_), .C(_15153_), .Y(_15154_) );
AOI21X1 AOI21X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_15150_), .B(_15154_), .C(_15015_), .Y(_15155_) );
INVX1 INVX1_2113 ( .gnd(gnd), .vdd(vdd), .A(_14536_), .Y(_15157_) );
AOI21X1 AOI21X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_14539_), .B(_14468_), .C(_15157_), .Y(_15158_) );
AOI21X1 AOI21X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_15152_), .B(_15153_), .C(_15151_), .Y(_15159_) );
AOI21X1 AOI21X1_2120 ( .gnd(gnd), .vdd(vdd), .A(_15144_), .B(_15149_), .C(_14537_), .Y(_15160_) );
NOR3X1 NOR3X1_445 ( .gnd(gnd), .vdd(vdd), .A(_15159_), .B(_15158_), .C(_15160_), .Y(_15161_) );
OAI21X1 OAI21X1_2408 ( .gnd(gnd), .vdd(vdd), .A(_15161_), .B(_15155_), .C(_15014_), .Y(_15162_) );
INVX1 INVX1_2114 ( .gnd(gnd), .vdd(vdd), .A(_15014_), .Y(_15163_) );
OAI21X1 OAI21X1_2409 ( .gnd(gnd), .vdd(vdd), .A(_15159_), .B(_15160_), .C(_15158_), .Y(_15164_) );
NAND3X1 NAND3X1_3410 ( .gnd(gnd), .vdd(vdd), .A(_15150_), .B(_15154_), .C(_15015_), .Y(_15165_) );
NAND3X1 NAND3X1_3411 ( .gnd(gnd), .vdd(vdd), .A(_15163_), .B(_15165_), .C(_15164_), .Y(_15166_) );
NAND3X1 NAND3X1_3412 ( .gnd(gnd), .vdd(vdd), .A(_15012_), .B(_15166_), .C(_15162_), .Y(_15168_) );
NAND3X1 NAND3X1_3413 ( .gnd(gnd), .vdd(vdd), .A(_15014_), .B(_15165_), .C(_15164_), .Y(_15169_) );
OAI21X1 OAI21X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_15161_), .B(_15155_), .C(_15163_), .Y(_15170_) );
NAND3X1 NAND3X1_3414 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf2_), .B(_15169_), .C(_15170_), .Y(_15171_) );
AOI21X1 AOI21X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15171_), .C(_15011_), .Y(_15172_) );
NAND3X1 NAND3X1_3415 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf1_), .B(_15166_), .C(_15162_), .Y(_15173_) );
NAND3X1 NAND3X1_3416 ( .gnd(gnd), .vdd(vdd), .A(_15012_), .B(_15169_), .C(_15170_), .Y(_15174_) );
AOI21X1 AOI21X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_15173_), .B(_15174_), .C(_14548_), .Y(_15175_) );
OAI21X1 OAI21X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .B(_15175_), .C(_15010_), .Y(_15176_) );
NAND2X1 NAND2X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_14547_), .B(_14551_), .Y(_15177_) );
NAND3X1 NAND3X1_3417 ( .gnd(gnd), .vdd(vdd), .A(_14548_), .B(_15173_), .C(_15174_), .Y(_15179_) );
NAND3X1 NAND3X1_3418 ( .gnd(gnd), .vdd(vdd), .A(_15011_), .B(_15168_), .C(_15171_), .Y(_15180_) );
NAND3X1 NAND3X1_3419 ( .gnd(gnd), .vdd(vdd), .A(_15177_), .B(_15179_), .C(_15180_), .Y(_15181_) );
NAND3X1 NAND3X1_3420 ( .gnd(gnd), .vdd(vdd), .A(_15485_), .B(_15181_), .C(_15176_), .Y(_15182_) );
AOI21X1 AOI21X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_15179_), .B(_15180_), .C(_15177_), .Y(_15183_) );
NOR3X1 NOR3X1_446 ( .gnd(gnd), .vdd(vdd), .A(_15175_), .B(_15010_), .C(_15172_), .Y(_15184_) );
OAI21X1 OAI21X1_2412 ( .gnd(gnd), .vdd(vdd), .A(_15184_), .B(_15183_), .C(_15101_), .Y(_15185_) );
NAND2X1 NAND2X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_15182_), .B(_15185_), .Y(_15186_) );
NAND3X1 NAND3X1_3421 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_140_), .B(_13207_), .C(_15186_), .Y(_15187_) );
INVX1 INVX1_2115 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_140_), .Y(_15188_) );
OAI21X1 OAI21X1_2413 ( .gnd(gnd), .vdd(vdd), .A(_15184_), .B(_15183_), .C(_15485_), .Y(_15190_) );
NAND3X1 NAND3X1_3422 ( .gnd(gnd), .vdd(vdd), .A(_15101_), .B(_15181_), .C(_15176_), .Y(_15191_) );
NAND3X1 NAND3X1_3423 ( .gnd(gnd), .vdd(vdd), .A(_13207_), .B(_15191_), .C(_15190_), .Y(_15192_) );
NAND2X1 NAND2X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_15188_), .B(_15192_), .Y(_15193_) );
AOI21X1 AOI21X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_15187_), .B(_15193_), .C(_15009_), .Y(_15194_) );
INVX1 INVX1_2116 ( .gnd(gnd), .vdd(vdd), .A(_15009_), .Y(_15195_) );
NAND2X1 NAND2X1_1976 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_140_), .B(_15192_), .Y(_15196_) );
NAND3X1 NAND3X1_3424 ( .gnd(gnd), .vdd(vdd), .A(_15188_), .B(_13207_), .C(_15186_), .Y(_15197_) );
AOI21X1 AOI21X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_15196_), .B(_15197_), .C(_15195_), .Y(_15198_) );
OAI21X1 OAI21X1_2414 ( .gnd(gnd), .vdd(vdd), .A(_15198_), .B(_15194_), .C(_15008_), .Y(_15199_) );
NAND3X1 NAND3X1_3425 ( .gnd(gnd), .vdd(vdd), .A(_15195_), .B(_15196_), .C(_15197_), .Y(_15201_) );
NAND3X1 NAND3X1_3426 ( .gnd(gnd), .vdd(vdd), .A(_15009_), .B(_15187_), .C(_15193_), .Y(_15202_) );
NAND3X1 NAND3X1_3427 ( .gnd(gnd), .vdd(vdd), .A(_15007_), .B(_15201_), .C(_15202_), .Y(_15203_) );
NAND3X1 NAND3X1_3428 ( .gnd(gnd), .vdd(vdd), .A(_15134_), .B(_15203_), .C(_15199_), .Y(_15204_) );
NAND2X1 NAND2X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_15203_), .B(_15199_), .Y(_15205_) );
AOI21X1 AOI21X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_15452_), .B(_15205_), .C(_13236_), .Y(_15206_) );
NAND3X1 NAND3X1_3429 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_156_), .B(_15204_), .C(_15206_), .Y(_15207_) );
INVX1 INVX1_2117 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_156_), .Y(_15208_) );
AOI21X1 AOI21X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_15201_), .B(_15202_), .C(_15007_), .Y(_15209_) );
NOR3X1 NOR3X1_447 ( .gnd(gnd), .vdd(vdd), .A(_15194_), .B(_15198_), .C(_15008_), .Y(_15210_) );
OAI21X1 OAI21X1_2415 ( .gnd(gnd), .vdd(vdd), .A(_15210_), .B(_15209_), .C(_15452_), .Y(_15212_) );
NAND3X1 NAND3X1_3430 ( .gnd(gnd), .vdd(vdd), .A(_13233_), .B(_15204_), .C(_15212_), .Y(_15213_) );
NAND2X1 NAND2X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_15208_), .B(_15213_), .Y(_15214_) );
AOI21X1 AOI21X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_15207_), .B(_15214_), .C(_14568_), .Y(_15215_) );
NAND2X1 NAND2X1_1979 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_156_), .B(_15213_), .Y(_15216_) );
NAND3X1 NAND3X1_3431 ( .gnd(gnd), .vdd(vdd), .A(_15208_), .B(_15204_), .C(_15206_), .Y(_15217_) );
AOI21X1 AOI21X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_15217_), .B(_15216_), .C(_14566_), .Y(_15218_) );
OAI21X1 OAI21X1_2416 ( .gnd(gnd), .vdd(vdd), .A(_15218_), .B(_15215_), .C(_15006_), .Y(_15219_) );
NAND3X1 NAND3X1_3432 ( .gnd(gnd), .vdd(vdd), .A(_14250_), .B(_14564_), .C(_14568_), .Y(_15220_) );
OAI21X1 OAI21X1_2417 ( .gnd(gnd), .vdd(vdd), .A(_14572_), .B(_14569_), .C(_15220_), .Y(_15221_) );
NAND3X1 NAND3X1_3433 ( .gnd(gnd), .vdd(vdd), .A(_14566_), .B(_15217_), .C(_15216_), .Y(_15223_) );
NAND3X1 NAND3X1_3434 ( .gnd(gnd), .vdd(vdd), .A(_14568_), .B(_15207_), .C(_15214_), .Y(_15224_) );
NAND3X1 NAND3X1_3435 ( .gnd(gnd), .vdd(vdd), .A(_15221_), .B(_15223_), .C(_15224_), .Y(_15225_) );
AOI21X1 AOI21X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_15225_), .B(_15219_), .C(_15167_), .Y(_15226_) );
NAND2X1 NAND2X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_15225_), .B(_15219_), .Y(_15227_) );
OAI21X1 OAI21X1_2418 ( .gnd(gnd), .vdd(vdd), .A(_15227_), .B(_15419_), .C(_13258_), .Y(_15228_) );
OAI21X1 OAI21X1_2419 ( .gnd(gnd), .vdd(vdd), .A(_15228_), .B(_15226_), .C(module_3_W_172_), .Y(_15229_) );
INVX1 INVX1_2118 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_172_), .Y(_15230_) );
NAND3X1 NAND3X1_3436 ( .gnd(gnd), .vdd(vdd), .A(_15419_), .B(_15225_), .C(_15219_), .Y(_15231_) );
AOI21X1 AOI21X1_2131 ( .gnd(gnd), .vdd(vdd), .A(_15223_), .B(_15224_), .C(_15221_), .Y(_15232_) );
NOR3X1 NOR3X1_448 ( .gnd(gnd), .vdd(vdd), .A(_15215_), .B(_15006_), .C(_15218_), .Y(_15234_) );
OAI21X1 OAI21X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_15234_), .B(_15232_), .C(_15167_), .Y(_15235_) );
NAND2X1 NAND2X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_15231_), .B(_15235_), .Y(_15236_) );
NAND3X1 NAND3X1_3437 ( .gnd(gnd), .vdd(vdd), .A(_15230_), .B(_13258_), .C(_15236_), .Y(_15237_) );
NAND3X1 NAND3X1_3438 ( .gnd(gnd), .vdd(vdd), .A(_15004_), .B(_15229_), .C(_15237_), .Y(_15238_) );
NAND3X1 NAND3X1_3439 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_172_), .B(_13258_), .C(_15236_), .Y(_15239_) );
OAI21X1 OAI21X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_15228_), .B(_15226_), .C(_15230_), .Y(_15240_) );
NAND3X1 NAND3X1_3440 ( .gnd(gnd), .vdd(vdd), .A(_14577_), .B(_15240_), .C(_15239_), .Y(_15241_) );
AOI21X1 AOI21X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_15238_), .B(_15241_), .C(_15003_), .Y(_15242_) );
INVX1 INVX1_2119 ( .gnd(gnd), .vdd(vdd), .A(_14580_), .Y(_15243_) );
AOI21X1 AOI21X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_15243_), .B(_14460_), .C(_14579_), .Y(_15245_) );
AOI21X1 AOI21X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_15240_), .B(_15239_), .C(_14577_), .Y(_15246_) );
AOI21X1 AOI21X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_15229_), .B(_15237_), .C(_15004_), .Y(_15247_) );
NOR3X1 NOR3X1_449 ( .gnd(gnd), .vdd(vdd), .A(_15246_), .B(_15247_), .C(_15245_), .Y(_15248_) );
OAI21X1 OAI21X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_15248_), .B(_15242_), .C(_15397_), .Y(_15249_) );
OAI21X1 OAI21X1_2423 ( .gnd(gnd), .vdd(vdd), .A(_15247_), .B(_15246_), .C(_15245_), .Y(_15250_) );
NAND3X1 NAND3X1_3441 ( .gnd(gnd), .vdd(vdd), .A(_15003_), .B(_15238_), .C(_15241_), .Y(_15251_) );
NAND3X1 NAND3X1_3442 ( .gnd(gnd), .vdd(vdd), .A(_15200_), .B(_15251_), .C(_15250_), .Y(_15252_) );
NAND3X1 NAND3X1_3443 ( .gnd(gnd), .vdd(vdd), .A(_13277_), .B(_15252_), .C(_15249_), .Y(_15253_) );
NAND2X1 NAND2X1_1982 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_188_), .B(_15253_), .Y(_15254_) );
INVX1 INVX1_2120 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_188_), .Y(_15256_) );
NAND3X1 NAND3X1_3444 ( .gnd(gnd), .vdd(vdd), .A(_15397_), .B(_15251_), .C(_15250_), .Y(_15257_) );
OAI21X1 OAI21X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_15248_), .B(_15242_), .C(_15200_), .Y(_15258_) );
NAND2X1 NAND2X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_15257_), .B(_15258_), .Y(_15259_) );
NAND3X1 NAND3X1_3445 ( .gnd(gnd), .vdd(vdd), .A(_15256_), .B(_13277_), .C(_15259_), .Y(_15260_) );
NAND3X1 NAND3X1_3446 ( .gnd(gnd), .vdd(vdd), .A(_15000_), .B(_15254_), .C(_15260_), .Y(_15261_) );
NAND3X1 NAND3X1_3447 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_188_), .B(_13277_), .C(_15259_), .Y(_15262_) );
NAND2X1 NAND2X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_15256_), .B(_15253_), .Y(_15263_) );
NAND3X1 NAND3X1_3448 ( .gnd(gnd), .vdd(vdd), .A(_14587_), .B(_15262_), .C(_15263_), .Y(_15264_) );
AOI21X1 AOI21X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_15261_), .B(_15264_), .C(_14999_), .Y(_15265_) );
INVX1 INVX1_2121 ( .gnd(gnd), .vdd(vdd), .A(_14590_), .Y(_15267_) );
AOI21X1 AOI21X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_14457_), .B(_15267_), .C(_14589_), .Y(_15268_) );
AOI21X1 AOI21X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_15262_), .B(_15263_), .C(_14587_), .Y(_15269_) );
AOI21X1 AOI21X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_15254_), .B(_15260_), .C(_15000_), .Y(_15270_) );
NOR3X1 NOR3X1_450 ( .gnd(gnd), .vdd(vdd), .A(_15269_), .B(_15270_), .C(_15268_), .Y(_15271_) );
OAI21X1 OAI21X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_15271_), .B(_15265_), .C(_15233_), .Y(_15272_) );
OAI21X1 OAI21X1_2426 ( .gnd(gnd), .vdd(vdd), .A(_15270_), .B(_15269_), .C(_15268_), .Y(_15273_) );
NAND3X1 NAND3X1_3449 ( .gnd(gnd), .vdd(vdd), .A(_14999_), .B(_15261_), .C(_15264_), .Y(_15274_) );
NAND3X1 NAND3X1_3450 ( .gnd(gnd), .vdd(vdd), .A(_15364_), .B(_15274_), .C(_15273_), .Y(_15275_) );
NAND2X1 NAND2X1_1985 ( .gnd(gnd), .vdd(vdd), .A(_15275_), .B(_15272_), .Y(_15276_) );
NAND3X1 NAND3X1_3451 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_204_), .B(_13304_), .C(_15276_), .Y(_15278_) );
INVX1 INVX1_2122 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_204_), .Y(_15279_) );
AOI21X1 AOI21X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_15274_), .B(_15273_), .C(_15233_), .Y(_15280_) );
NAND2X1 NAND2X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_15274_), .B(_15273_), .Y(_15281_) );
OAI21X1 OAI21X1_2427 ( .gnd(gnd), .vdd(vdd), .A(_15281_), .B(_15364_), .C(_13304_), .Y(_15282_) );
OAI21X1 OAI21X1_2428 ( .gnd(gnd), .vdd(vdd), .A(_15282_), .B(_15280_), .C(_15279_), .Y(_15283_) );
AOI21X1 AOI21X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_15283_), .B(_15278_), .C(_14598_), .Y(_15284_) );
OAI21X1 OAI21X1_2429 ( .gnd(gnd), .vdd(vdd), .A(_15282_), .B(_15280_), .C(module_3_W_204_), .Y(_15285_) );
NAND3X1 NAND3X1_3452 ( .gnd(gnd), .vdd(vdd), .A(_15279_), .B(_13304_), .C(_15276_), .Y(_15286_) );
AOI21X1 AOI21X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_15285_), .B(_15286_), .C(_14597_), .Y(_15287_) );
OAI21X1 OAI21X1_2430 ( .gnd(gnd), .vdd(vdd), .A(_15287_), .B(_15284_), .C(_14998_), .Y(_15289_) );
AOI21X1 AOI21X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_14596_), .B(_14598_), .C(_14360_), .Y(_15290_) );
OAI21X1 OAI21X1_2431 ( .gnd(gnd), .vdd(vdd), .A(_15290_), .B(_14455_), .C(_14599_), .Y(_15291_) );
NAND3X1 NAND3X1_3453 ( .gnd(gnd), .vdd(vdd), .A(_14597_), .B(_15285_), .C(_15286_), .Y(_15292_) );
NAND3X1 NAND3X1_3454 ( .gnd(gnd), .vdd(vdd), .A(_14598_), .B(_15283_), .C(_15278_), .Y(_15293_) );
NAND3X1 NAND3X1_3455 ( .gnd(gnd), .vdd(vdd), .A(_15292_), .B(_15293_), .C(_15291_), .Y(_15294_) );
NAND3X1 NAND3X1_3456 ( .gnd(gnd), .vdd(vdd), .A(_15343_), .B(_15294_), .C(_15289_), .Y(_15295_) );
AOI21X1 AOI21X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_15292_), .B(_15293_), .C(_15291_), .Y(_15296_) );
NOR3X1 NOR3X1_451 ( .gnd(gnd), .vdd(vdd), .A(_15284_), .B(_14998_), .C(_15287_), .Y(_15297_) );
OAI21X1 OAI21X1_2432 ( .gnd(gnd), .vdd(vdd), .A(_15297_), .B(_15296_), .C(_15266_), .Y(_15298_) );
NAND2X1 NAND2X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_15295_), .B(_15298_), .Y(_15300_) );
NAND3X1 NAND3X1_3457 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_220_), .B(_13325_), .C(_15300_), .Y(_15301_) );
INVX1 INVX1_2123 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_220_), .Y(_15302_) );
AOI21X1 AOI21X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_15294_), .B(_15289_), .C(_15266_), .Y(_15303_) );
NAND2X1 NAND2X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_15294_), .B(_15289_), .Y(_15304_) );
OAI21X1 OAI21X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_15304_), .B(_15343_), .C(_13325_), .Y(_15305_) );
OAI21X1 OAI21X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_15305_), .B(_15303_), .C(_15302_), .Y(_15306_) );
AOI21X1 AOI21X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_15306_), .B(_15301_), .C(_14611_), .Y(_15307_) );
OAI21X1 OAI21X1_2435 ( .gnd(gnd), .vdd(vdd), .A(_15305_), .B(_15303_), .C(module_3_W_220_), .Y(_15308_) );
NAND3X1 NAND3X1_3458 ( .gnd(gnd), .vdd(vdd), .A(_15302_), .B(_13325_), .C(_15300_), .Y(_15309_) );
AOI21X1 AOI21X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_15308_), .B(_15309_), .C(_14608_), .Y(_15311_) );
OAI21X1 OAI21X1_2436 ( .gnd(gnd), .vdd(vdd), .A(_15307_), .B(_15311_), .C(_14996_), .Y(_15312_) );
AOI21X1 AOI21X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_14394_), .B(_14402_), .C(_14404_), .Y(_15313_) );
NAND3X1 NAND3X1_3459 ( .gnd(gnd), .vdd(vdd), .A(_14397_), .B(_14611_), .C(_14610_), .Y(_15314_) );
OAI21X1 OAI21X1_2437 ( .gnd(gnd), .vdd(vdd), .A(_15313_), .B(_14612_), .C(_15314_), .Y(_15315_) );
NAND3X1 NAND3X1_3460 ( .gnd(gnd), .vdd(vdd), .A(_14608_), .B(_15308_), .C(_15309_), .Y(_15316_) );
NAND3X1 NAND3X1_3461 ( .gnd(gnd), .vdd(vdd), .A(_14611_), .B(_15306_), .C(_15301_), .Y(_15317_) );
NAND3X1 NAND3X1_3462 ( .gnd(gnd), .vdd(vdd), .A(_15315_), .B(_15316_), .C(_15317_), .Y(_15318_) );
AOI21X1 AOI21X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_15318_), .B(_15312_), .C(_15299_), .Y(_15319_) );
NAND2X1 NAND2X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_15318_), .B(_15312_), .Y(_15320_) );
OAI21X1 OAI21X1_2438 ( .gnd(gnd), .vdd(vdd), .A(_15320_), .B(_15310_), .C(_13351_), .Y(_15322_) );
OAI21X1 OAI21X1_2439 ( .gnd(gnd), .vdd(vdd), .A(_15322_), .B(_15319_), .C(module_3_W_236_), .Y(_15323_) );
INVX1 INVX1_2124 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_236_), .Y(_15324_) );
NAND3X1 NAND3X1_3463 ( .gnd(gnd), .vdd(vdd), .A(_15310_), .B(_15318_), .C(_15312_), .Y(_15325_) );
AOI21X1 AOI21X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_15316_), .B(_15317_), .C(_15315_), .Y(_15326_) );
NOR3X1 NOR3X1_452 ( .gnd(gnd), .vdd(vdd), .A(_15307_), .B(_14996_), .C(_15311_), .Y(_15327_) );
OAI21X1 OAI21X1_2440 ( .gnd(gnd), .vdd(vdd), .A(_15327_), .B(_15326_), .C(_15299_), .Y(_15328_) );
NAND2X1 NAND2X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_15325_), .B(_15328_), .Y(_15329_) );
NAND3X1 NAND3X1_3464 ( .gnd(gnd), .vdd(vdd), .A(_15324_), .B(_13351_), .C(_15329_), .Y(_15330_) );
NAND3X1 NAND3X1_3465 ( .gnd(gnd), .vdd(vdd), .A(_14994_), .B(_15323_), .C(_15330_), .Y(_15331_) );
NAND3X1 NAND3X1_3466 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_236_), .B(_13351_), .C(_15329_), .Y(_15333_) );
OAI21X1 OAI21X1_2441 ( .gnd(gnd), .vdd(vdd), .A(_15322_), .B(_15319_), .C(_15324_), .Y(_15334_) );
NAND3X1 NAND3X1_3467 ( .gnd(gnd), .vdd(vdd), .A(_14618_), .B(_15334_), .C(_15333_), .Y(_15335_) );
AOI21X1 AOI21X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_15331_), .B(_15335_), .C(_14993_), .Y(_15336_) );
INVX1 INVX1_2125 ( .gnd(gnd), .vdd(vdd), .A(_14621_), .Y(_15337_) );
AOI21X1 AOI21X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_14624_), .B(_15337_), .C(_14620_), .Y(_15338_) );
NAND3X1 NAND3X1_3468 ( .gnd(gnd), .vdd(vdd), .A(_14994_), .B(_15334_), .C(_15333_), .Y(_15339_) );
NAND3X1 NAND3X1_3469 ( .gnd(gnd), .vdd(vdd), .A(_14618_), .B(_15323_), .C(_15330_), .Y(_15340_) );
AOI21X1 AOI21X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_15339_), .B(_15340_), .C(_15338_), .Y(_15341_) );
OAI21X1 OAI21X1_2442 ( .gnd(gnd), .vdd(vdd), .A(_15341_), .B(_15336_), .C(_16544_), .Y(_15342_) );
AOI21X1 AOI21X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_15334_), .B(_15333_), .C(_14618_), .Y(_15344_) );
AOI21X1 AOI21X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_15323_), .B(_15330_), .C(_14994_), .Y(_15345_) );
OAI21X1 OAI21X1_2443 ( .gnd(gnd), .vdd(vdd), .A(_15344_), .B(_15345_), .C(_15338_), .Y(_15346_) );
NAND3X1 NAND3X1_3470 ( .gnd(gnd), .vdd(vdd), .A(_14993_), .B(_15331_), .C(_15335_), .Y(_15347_) );
NAND3X1 NAND3X1_3471 ( .gnd(gnd), .vdd(vdd), .A(_16545_), .B(_15347_), .C(_15346_), .Y(_15348_) );
NAND2X1 NAND2X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_15348_), .B(_15342_), .Y(_15349_) );
NAND3X1 NAND3X1_3472 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_252_), .B(_13375_), .C(_15349_), .Y(_15350_) );
INVX1 INVX1_2126 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_252_), .Y(_15351_) );
AOI21X1 AOI21X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_15347_), .B(_15346_), .C(_16544_), .Y(_15352_) );
NAND2X1 NAND2X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_15347_), .B(_15346_), .Y(_15353_) );
OAI21X1 OAI21X1_2444 ( .gnd(gnd), .vdd(vdd), .A(_15353_), .B(_16545_), .C(_13375_), .Y(_15355_) );
OAI21X1 OAI21X1_2445 ( .gnd(gnd), .vdd(vdd), .A(_15355_), .B(_15352_), .C(_15351_), .Y(_15356_) );
AOI21X1 AOI21X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_15356_), .B(_15350_), .C(_14985_), .Y(_15357_) );
INVX1 INVX1_2127 ( .gnd(gnd), .vdd(vdd), .A(_15357_), .Y(_15358_) );
NAND3X1 NAND3X1_3473 ( .gnd(gnd), .vdd(vdd), .A(_14985_), .B(_15356_), .C(_15350_), .Y(_15359_) );
NAND2X1 NAND2X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_15359_), .B(_15358_), .Y(_15360_) );
XOR2X1 XOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_15360_), .B(_14992_), .Y(module_3_H_20_) );
OAI21X1 OAI21X1_2446 ( .gnd(gnd), .vdd(vdd), .A(_15357_), .B(_14992_), .C(_15359_), .Y(_15361_) );
NAND2X1 NAND2X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_13375_), .B(_15349_), .Y(_15362_) );
NOR2X1 NOR2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_252_), .B(_15362_), .Y(_15363_) );
AOI21X1 AOI21X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_14993_), .B(_15335_), .C(_15344_), .Y(_15365_) );
INVX1 INVX1_2128 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_237_), .Y(_15366_) );
OAI21X1 OAI21X1_2447 ( .gnd(gnd), .vdd(vdd), .A(_15311_), .B(_14996_), .C(_15316_), .Y(_15367_) );
INVX1 INVX1_2129 ( .gnd(gnd), .vdd(vdd), .A(_15308_), .Y(_15368_) );
AOI21X1 AOI21X1_2159 ( .gnd(gnd), .vdd(vdd), .A(_15293_), .B(_15291_), .C(_15284_), .Y(_15369_) );
INVX1 INVX1_2130 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_205_), .Y(_15370_) );
OAI21X1 OAI21X1_2448 ( .gnd(gnd), .vdd(vdd), .A(_15268_), .B(_15270_), .C(_15261_), .Y(_15371_) );
INVX1 INVX1_2131 ( .gnd(gnd), .vdd(vdd), .A(_15254_), .Y(_15372_) );
AOI21X1 AOI21X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_15003_), .B(_15241_), .C(_15246_), .Y(_15373_) );
INVX1 INVX1_2132 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_173_), .Y(_15374_) );
INVX1 INVX1_2133 ( .gnd(gnd), .vdd(vdd), .A(_16315_), .Y(_15376_) );
AOI21X1 AOI21X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_15221_), .B(_15224_), .C(_15215_), .Y(_15377_) );
INVX1 INVX1_2134 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_157_), .Y(_15378_) );
INVX1 INVX1_2135 ( .gnd(gnd), .vdd(vdd), .A(_16231_), .Y(_15379_) );
AOI21X1 AOI21X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_15007_), .B(_15202_), .C(_15194_), .Y(_15380_) );
INVX1 INVX1_2136 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_141_), .Y(_15381_) );
OAI21X1 OAI21X1_2449 ( .gnd(gnd), .vdd(vdd), .A(_15175_), .B(_15010_), .C(_15179_), .Y(_15382_) );
INVX1 INVX1_2137 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf3_), .Y(_15383_) );
AOI21X1 AOI21X1_2163 ( .gnd(gnd), .vdd(vdd), .A(_15154_), .B(_15015_), .C(_15159_), .Y(_15384_) );
INVX1 INVX1_2138 ( .gnd(gnd), .vdd(vdd), .A(_15152_), .Y(_15385_) );
INVX1 INVX1_2139 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf1_), .Y(_15387_) );
AOI21X1 AOI21X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_15131_), .B(_15019_), .C(_15136_), .Y(_15388_) );
INVX1 INVX1_2140 ( .gnd(gnd), .vdd(vdd), .A(_15129_), .Y(_15389_) );
INVX1 INVX1_2141 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf1_), .Y(_15390_) );
AOI21X1 AOI21X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_15114_), .B(_15111_), .C(_15105_), .Y(_15391_) );
INVX1 INVX1_2142 ( .gnd(gnd), .vdd(vdd), .A(_15100_), .Y(_15392_) );
INVX1 INVX1_2143 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf1_), .Y(_15393_) );
OAI21X1 OAI21X1_2450 ( .gnd(gnd), .vdd(vdd), .A(_15026_), .B(_15087_), .C(_15091_), .Y(_15394_) );
INVX1 INVX1_2144 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf3_), .Y(_15395_) );
AOI21X1 AOI21X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_15066_), .B(_15031_), .C(_15071_), .Y(_15396_) );
INVX1 INVX1_2145 ( .gnd(gnd), .vdd(vdd), .A(_15064_), .Y(_15398_) );
INVX1 INVX1_2146 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf3_), .Y(_15399_) );
OAI21X1 OAI21X1_2451 ( .gnd(gnd), .vdd(vdd), .A(_15050_), .B(_15049_), .C(_15045_), .Y(_15400_) );
INVX1 INVX1_2147 ( .gnd(gnd), .vdd(vdd), .A(_15040_), .Y(_15401_) );
XOR2X1 XOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_12_), .B(module_3_W_13_), .Y(_15402_) );
INVX1 INVX1_2148 ( .gnd(gnd), .vdd(vdd), .A(_15402_), .Y(_15403_) );
OAI21X1 OAI21X1_2452 ( .gnd(gnd), .vdd(vdd), .A(_15683_), .B(_15694_), .C(module_3_W_9_), .Y(_15404_) );
NAND2X1 NAND2X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_13401_), .B(_13544_), .Y(_15405_) );
NAND2X1 NAND2X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_15404_), .B(_15405_), .Y(_15406_) );
NAND2X1 NAND2X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15406_), .Y(_15407_) );
NAND3X1 NAND3X1_3474 ( .gnd(gnd), .vdd(vdd), .A(_15402_), .B(_15404_), .C(_15405_), .Y(_15409_) );
AOI21X1 AOI21X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_15409_), .B(_15407_), .C(module_3_W_29_), .Y(_15410_) );
INVX1 INVX1_2149 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_29_), .Y(_15411_) );
NAND2X1 NAND2X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_15402_), .B(_15406_), .Y(_15412_) );
NAND3X1 NAND3X1_3475 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15404_), .C(_15405_), .Y(_15413_) );
AOI21X1 AOI21X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_15413_), .B(_15412_), .C(_15411_), .Y(_15414_) );
OAI21X1 OAI21X1_2453 ( .gnd(gnd), .vdd(vdd), .A(_15414_), .B(_15410_), .C(_15401_), .Y(_15415_) );
NAND3X1 NAND3X1_3476 ( .gnd(gnd), .vdd(vdd), .A(_15411_), .B(_15413_), .C(_15412_), .Y(_15416_) );
NAND3X1 NAND3X1_3477 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_29_), .B(_15409_), .C(_15407_), .Y(_15417_) );
NAND3X1 NAND3X1_3478 ( .gnd(gnd), .vdd(vdd), .A(_15040_), .B(_15417_), .C(_15416_), .Y(_15418_) );
NAND3X1 NAND3X1_3479 ( .gnd(gnd), .vdd(vdd), .A(_15415_), .B(_15418_), .C(_15400_), .Y(_15420_) );
AOI21X1 AOI21X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_15043_), .B(_15036_), .C(_15044_), .Y(_15421_) );
AOI21X1 AOI21X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_15417_), .B(_15416_), .C(_15040_), .Y(_15422_) );
NOR3X1 NOR3X1_453 ( .gnd(gnd), .vdd(vdd), .A(_15410_), .B(_15401_), .C(_15414_), .Y(_15423_) );
OAI21X1 OAI21X1_2454 ( .gnd(gnd), .vdd(vdd), .A(_15423_), .B(_15422_), .C(_15421_), .Y(_15424_) );
XNOR2X1 XNOR2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_13407_), .B(_15770_), .Y(_15425_) );
INVX1 INVX1_2150 ( .gnd(gnd), .vdd(vdd), .A(_15425_), .Y(_15426_) );
NAND3X1 NAND3X1_3480 ( .gnd(gnd), .vdd(vdd), .A(_15424_), .B(_15426_), .C(_15420_), .Y(_15427_) );
NOR3X1 NOR3X1_454 ( .gnd(gnd), .vdd(vdd), .A(_15421_), .B(_15422_), .C(_15423_), .Y(_15428_) );
AOI21X1 AOI21X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_15415_), .B(_15418_), .C(_15400_), .Y(_15429_) );
OAI21X1 OAI21X1_2455 ( .gnd(gnd), .vdd(vdd), .A(_15428_), .B(_15429_), .C(_15425_), .Y(_15431_) );
NAND3X1 NAND3X1_3481 ( .gnd(gnd), .vdd(vdd), .A(_15399_), .B(_15427_), .C(_15431_), .Y(_15432_) );
NAND3X1 NAND3X1_3482 ( .gnd(gnd), .vdd(vdd), .A(_15424_), .B(_15425_), .C(_15420_), .Y(_15433_) );
OAI21X1 OAI21X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_15428_), .B(_15429_), .C(_15426_), .Y(_15434_) );
NAND3X1 NAND3X1_3483 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf2_), .B(_15433_), .C(_15434_), .Y(_15435_) );
NAND3X1 NAND3X1_3484 ( .gnd(gnd), .vdd(vdd), .A(_15398_), .B(_15432_), .C(_15435_), .Y(_15436_) );
AOI21X1 AOI21X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_15433_), .B(_15434_), .C(bloque_datos_13_bF_buf1_), .Y(_15437_) );
AOI21X1 AOI21X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_15427_), .B(_15431_), .C(_15399_), .Y(_15438_) );
OAI21X1 OAI21X1_2457 ( .gnd(gnd), .vdd(vdd), .A(_15437_), .B(_15438_), .C(_15064_), .Y(_15439_) );
NAND3X1 NAND3X1_3485 ( .gnd(gnd), .vdd(vdd), .A(_15436_), .B(_15439_), .C(_15396_), .Y(_15440_) );
OAI21X1 OAI21X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_15072_), .B(_15070_), .C(_15062_), .Y(_15442_) );
NAND3X1 NAND3X1_3486 ( .gnd(gnd), .vdd(vdd), .A(_15064_), .B(_15432_), .C(_15435_), .Y(_15443_) );
OAI21X1 OAI21X1_2459 ( .gnd(gnd), .vdd(vdd), .A(_15437_), .B(_15438_), .C(_15398_), .Y(_15444_) );
NAND3X1 NAND3X1_3487 ( .gnd(gnd), .vdd(vdd), .A(_15443_), .B(_15444_), .C(_15442_), .Y(_15445_) );
XNOR2X1 XNOR2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_13607_), .B(_15814_), .Y(_15446_) );
INVX1 INVX1_2151 ( .gnd(gnd), .vdd(vdd), .A(_15446_), .Y(_15447_) );
NAND3X1 NAND3X1_3488 ( .gnd(gnd), .vdd(vdd), .A(_15445_), .B(_15447_), .C(_15440_), .Y(_15448_) );
AOI21X1 AOI21X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_15443_), .B(_15444_), .C(_15442_), .Y(_15449_) );
AOI21X1 AOI21X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_15436_), .B(_15439_), .C(_15396_), .Y(_15450_) );
OAI21X1 OAI21X1_2460 ( .gnd(gnd), .vdd(vdd), .A(_15450_), .B(_15449_), .C(_15446_), .Y(_15451_) );
NAND3X1 NAND3X1_3489 ( .gnd(gnd), .vdd(vdd), .A(_15395_), .B(_15448_), .C(_15451_), .Y(_15453_) );
NOR3X1 NOR3X1_455 ( .gnd(gnd), .vdd(vdd), .A(_15449_), .B(_15446_), .C(_15450_), .Y(_15454_) );
AOI21X1 AOI21X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_15445_), .B(_15440_), .C(_15447_), .Y(_15455_) );
OAI21X1 OAI21X1_2461 ( .gnd(gnd), .vdd(vdd), .A(_15454_), .B(_15455_), .C(bloque_datos_29_bF_buf2_), .Y(_15456_) );
NAND3X1 NAND3X1_3490 ( .gnd(gnd), .vdd(vdd), .A(_15078_), .B(_15453_), .C(_15456_), .Y(_15457_) );
INVX1 INVX1_2152 ( .gnd(gnd), .vdd(vdd), .A(_15078_), .Y(_15458_) );
NOR3X1 NOR3X1_456 ( .gnd(gnd), .vdd(vdd), .A(_15455_), .B(bloque_datos_29_bF_buf1_), .C(_15454_), .Y(_15459_) );
AOI21X1 AOI21X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_15448_), .B(_15451_), .C(_15395_), .Y(_15460_) );
OAI21X1 OAI21X1_2462 ( .gnd(gnd), .vdd(vdd), .A(_15459_), .B(_15460_), .C(_15458_), .Y(_15461_) );
AOI21X1 AOI21X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_15457_), .B(_15461_), .C(_15394_), .Y(_15462_) );
AOI21X1 AOI21X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_15092_), .B(_15089_), .C(_15083_), .Y(_15464_) );
NAND3X1 NAND3X1_3491 ( .gnd(gnd), .vdd(vdd), .A(_15458_), .B(_15453_), .C(_15456_), .Y(_15465_) );
OAI21X1 OAI21X1_2463 ( .gnd(gnd), .vdd(vdd), .A(_15459_), .B(_15460_), .C(_15078_), .Y(_15466_) );
AOI21X1 AOI21X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_15465_), .B(_15466_), .C(_15464_), .Y(_15467_) );
XNOR2X1 XNOR2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_13424_), .B(_15869_), .Y(_15468_) );
NOR3X1 NOR3X1_457 ( .gnd(gnd), .vdd(vdd), .A(_15467_), .B(_15468_), .C(_15462_), .Y(_15469_) );
NAND3X1 NAND3X1_3492 ( .gnd(gnd), .vdd(vdd), .A(_15465_), .B(_15464_), .C(_15466_), .Y(_15470_) );
NAND3X1 NAND3X1_3493 ( .gnd(gnd), .vdd(vdd), .A(_15394_), .B(_15457_), .C(_15461_), .Y(_15471_) );
INVX1 INVX1_2153 ( .gnd(gnd), .vdd(vdd), .A(_15468_), .Y(_15472_) );
AOI21X1 AOI21X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_15470_), .B(_15471_), .C(_15472_), .Y(_15473_) );
OAI21X1 OAI21X1_2464 ( .gnd(gnd), .vdd(vdd), .A(_15469_), .B(_15473_), .C(_15393_), .Y(_15475_) );
NAND3X1 NAND3X1_3494 ( .gnd(gnd), .vdd(vdd), .A(_15472_), .B(_15470_), .C(_15471_), .Y(_15476_) );
OAI21X1 OAI21X1_2465 ( .gnd(gnd), .vdd(vdd), .A(_15462_), .B(_15467_), .C(_15468_), .Y(_15477_) );
NAND3X1 NAND3X1_3495 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf0_), .B(_15476_), .C(_15477_), .Y(_15478_) );
NAND3X1 NAND3X1_3496 ( .gnd(gnd), .vdd(vdd), .A(_15392_), .B(_15478_), .C(_15475_), .Y(_15479_) );
AOI21X1 AOI21X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_15476_), .B(_15477_), .C(bloque_datos_45_bF_buf4_), .Y(_15480_) );
NOR3X1 NOR3X1_458 ( .gnd(gnd), .vdd(vdd), .A(_15473_), .B(_15393_), .C(_15469_), .Y(_15481_) );
OAI21X1 OAI21X1_2466 ( .gnd(gnd), .vdd(vdd), .A(_15481_), .B(_15480_), .C(_15100_), .Y(_15482_) );
NAND3X1 NAND3X1_3497 ( .gnd(gnd), .vdd(vdd), .A(_15479_), .B(_15482_), .C(_15391_), .Y(_15483_) );
OAI21X1 OAI21X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_15022_), .B(_15108_), .C(_15113_), .Y(_15484_) );
NAND3X1 NAND3X1_3498 ( .gnd(gnd), .vdd(vdd), .A(_15100_), .B(_15478_), .C(_15475_), .Y(_15486_) );
OAI21X1 OAI21X1_2468 ( .gnd(gnd), .vdd(vdd), .A(_15481_), .B(_15480_), .C(_15392_), .Y(_15487_) );
NAND3X1 NAND3X1_3499 ( .gnd(gnd), .vdd(vdd), .A(_15486_), .B(_15484_), .C(_15487_), .Y(_15488_) );
XOR2X1 XOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_13432_), .B(_15946_), .Y(_15489_) );
INVX1 INVX1_2154 ( .gnd(gnd), .vdd(vdd), .A(_15489_), .Y(_15490_) );
NAND3X1 NAND3X1_3500 ( .gnd(gnd), .vdd(vdd), .A(_15490_), .B(_15488_), .C(_15483_), .Y(_15491_) );
AOI21X1 AOI21X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_15486_), .B(_15487_), .C(_15484_), .Y(_15492_) );
AOI21X1 AOI21X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_15479_), .B(_15482_), .C(_15391_), .Y(_15493_) );
OAI21X1 OAI21X1_2469 ( .gnd(gnd), .vdd(vdd), .A(_15493_), .B(_15492_), .C(_15489_), .Y(_15494_) );
NAND3X1 NAND3X1_3501 ( .gnd(gnd), .vdd(vdd), .A(_15390_), .B(_15491_), .C(_15494_), .Y(_15495_) );
NAND3X1 NAND3X1_3502 ( .gnd(gnd), .vdd(vdd), .A(_15489_), .B(_15488_), .C(_15483_), .Y(_15497_) );
OAI21X1 OAI21X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_15493_), .B(_15492_), .C(_15490_), .Y(_15498_) );
NAND3X1 NAND3X1_3503 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf0_), .B(_15497_), .C(_15498_), .Y(_15499_) );
NAND3X1 NAND3X1_3504 ( .gnd(gnd), .vdd(vdd), .A(_15389_), .B(_15495_), .C(_15499_), .Y(_15500_) );
AOI21X1 AOI21X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_15497_), .B(_15498_), .C(bloque_datos_61_bF_buf4_), .Y(_15501_) );
AOI21X1 AOI21X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_15491_), .B(_15494_), .C(_15390_), .Y(_15502_) );
OAI21X1 OAI21X1_2471 ( .gnd(gnd), .vdd(vdd), .A(_15501_), .B(_15502_), .C(_15129_), .Y(_15503_) );
NAND3X1 NAND3X1_3505 ( .gnd(gnd), .vdd(vdd), .A(_15500_), .B(_15503_), .C(_15388_), .Y(_15504_) );
OAI21X1 OAI21X1_2472 ( .gnd(gnd), .vdd(vdd), .A(_15135_), .B(_15137_), .C(_15127_), .Y(_15505_) );
NAND3X1 NAND3X1_3506 ( .gnd(gnd), .vdd(vdd), .A(_15129_), .B(_15495_), .C(_15499_), .Y(_15506_) );
OAI21X1 OAI21X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_15501_), .B(_15502_), .C(_15389_), .Y(_15508_) );
NAND3X1 NAND3X1_3507 ( .gnd(gnd), .vdd(vdd), .A(_15506_), .B(_15505_), .C(_15508_), .Y(_15509_) );
XNOR2X1 XNOR2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_13437_), .B(_16012_), .Y(_15510_) );
INVX1 INVX1_2155 ( .gnd(gnd), .vdd(vdd), .A(_15510_), .Y(_15511_) );
NAND3X1 NAND3X1_3508 ( .gnd(gnd), .vdd(vdd), .A(_15511_), .B(_15509_), .C(_15504_), .Y(_15512_) );
AOI21X1 AOI21X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_15506_), .B(_15508_), .C(_15505_), .Y(_15513_) );
AOI21X1 AOI21X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_15500_), .B(_15503_), .C(_15388_), .Y(_15514_) );
OAI21X1 OAI21X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_15513_), .B(_15514_), .C(_15510_), .Y(_15515_) );
NAND3X1 NAND3X1_3509 ( .gnd(gnd), .vdd(vdd), .A(_15387_), .B(_15512_), .C(_15515_), .Y(_15516_) );
NAND3X1 NAND3X1_3510 ( .gnd(gnd), .vdd(vdd), .A(_15510_), .B(_15509_), .C(_15504_), .Y(_15517_) );
OAI21X1 OAI21X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_15513_), .B(_15514_), .C(_15511_), .Y(_15519_) );
NAND3X1 NAND3X1_3511 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf0_), .B(_15517_), .C(_15519_), .Y(_15520_) );
NAND3X1 NAND3X1_3512 ( .gnd(gnd), .vdd(vdd), .A(_15385_), .B(_15516_), .C(_15520_), .Y(_15521_) );
AOI21X1 AOI21X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_15517_), .B(_15519_), .C(bloque_datos_77_bF_buf4_), .Y(_15522_) );
AOI21X1 AOI21X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_15512_), .B(_15515_), .C(_15387_), .Y(_15523_) );
OAI21X1 OAI21X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_15522_), .B(_15523_), .C(_15152_), .Y(_15524_) );
NAND3X1 NAND3X1_3513 ( .gnd(gnd), .vdd(vdd), .A(_15521_), .B(_15524_), .C(_15384_), .Y(_15525_) );
OAI21X1 OAI21X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_15160_), .B(_15158_), .C(_15150_), .Y(_15526_) );
NAND3X1 NAND3X1_3514 ( .gnd(gnd), .vdd(vdd), .A(_15152_), .B(_15516_), .C(_15520_), .Y(_15527_) );
OAI21X1 OAI21X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_15522_), .B(_15523_), .C(_15385_), .Y(_15528_) );
NAND3X1 NAND3X1_3515 ( .gnd(gnd), .vdd(vdd), .A(_15527_), .B(_15526_), .C(_15528_), .Y(_15530_) );
XNOR2X1 XNOR2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_13443_), .B(_16056_), .Y(_15531_) );
INVX1 INVX1_2156 ( .gnd(gnd), .vdd(vdd), .A(_15531_), .Y(_15532_) );
NAND3X1 NAND3X1_3516 ( .gnd(gnd), .vdd(vdd), .A(_15532_), .B(_15530_), .C(_15525_), .Y(_15533_) );
AOI21X1 AOI21X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_15527_), .B(_15528_), .C(_15526_), .Y(_15534_) );
AOI21X1 AOI21X1_2192 ( .gnd(gnd), .vdd(vdd), .A(_15521_), .B(_15524_), .C(_15384_), .Y(_15535_) );
OAI21X1 OAI21X1_2479 ( .gnd(gnd), .vdd(vdd), .A(_15534_), .B(_15535_), .C(_15531_), .Y(_15536_) );
NAND3X1 NAND3X1_3517 ( .gnd(gnd), .vdd(vdd), .A(_15383_), .B(_15533_), .C(_15536_), .Y(_15537_) );
NOR3X1 NOR3X1_459 ( .gnd(gnd), .vdd(vdd), .A(_15534_), .B(_15531_), .C(_15535_), .Y(_15538_) );
AOI21X1 AOI21X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_15530_), .B(_15525_), .C(_15532_), .Y(_15539_) );
OAI21X1 OAI21X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_15538_), .B(_15539_), .C(bloque_datos_93_bF_buf2_), .Y(_15541_) );
NAND3X1 NAND3X1_3518 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15537_), .C(_15541_), .Y(_15542_) );
INVX1 INVX1_2157 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .Y(_15543_) );
NOR3X1 NOR3X1_460 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf1_), .B(_15539_), .C(_15538_), .Y(_15544_) );
AOI21X1 AOI21X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_15533_), .B(_15536_), .C(_15383_), .Y(_15545_) );
OAI21X1 OAI21X1_2481 ( .gnd(gnd), .vdd(vdd), .A(_15544_), .B(_15545_), .C(_15543_), .Y(_15546_) );
AOI21X1 AOI21X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_15542_), .B(_15546_), .C(_15382_), .Y(_15547_) );
AOI21X1 AOI21X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_15177_), .B(_15180_), .C(_15172_), .Y(_15548_) );
NAND3X1 NAND3X1_3519 ( .gnd(gnd), .vdd(vdd), .A(_15543_), .B(_15537_), .C(_15541_), .Y(_15549_) );
OAI21X1 OAI21X1_2482 ( .gnd(gnd), .vdd(vdd), .A(_15544_), .B(_15545_), .C(_15168_), .Y(_15550_) );
AOI21X1 AOI21X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_15549_), .B(_15550_), .C(_15548_), .Y(_15552_) );
OAI21X1 OAI21X1_2483 ( .gnd(gnd), .vdd(vdd), .A(_15547_), .B(_15552_), .C(_16154_), .Y(_15553_) );
NAND3X1 NAND3X1_3520 ( .gnd(gnd), .vdd(vdd), .A(_15548_), .B(_15549_), .C(_15550_), .Y(_15554_) );
NAND3X1 NAND3X1_3521 ( .gnd(gnd), .vdd(vdd), .A(_15382_), .B(_15542_), .C(_15546_), .Y(_15555_) );
NAND3X1 NAND3X1_3522 ( .gnd(gnd), .vdd(vdd), .A(_16165_), .B(_15554_), .C(_15555_), .Y(_15556_) );
NAND2X1 NAND2X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_15556_), .B(_15553_), .Y(_15557_) );
NAND3X1 NAND3X1_3523 ( .gnd(gnd), .vdd(vdd), .A(_15381_), .B(_13450_), .C(_15557_), .Y(_15558_) );
OAI21X1 OAI21X1_2484 ( .gnd(gnd), .vdd(vdd), .A(_15547_), .B(_15552_), .C(_16165_), .Y(_15559_) );
NAND3X1 NAND3X1_3524 ( .gnd(gnd), .vdd(vdd), .A(_16154_), .B(_15554_), .C(_15555_), .Y(_15560_) );
NAND3X1 NAND3X1_3525 ( .gnd(gnd), .vdd(vdd), .A(_13450_), .B(_15560_), .C(_15559_), .Y(_15561_) );
NAND2X1 NAND2X1_2000 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_141_), .B(_15561_), .Y(_15563_) );
AOI21X1 AOI21X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_15558_), .B(_15563_), .C(_15196_), .Y(_15564_) );
INVX1 INVX1_2158 ( .gnd(gnd), .vdd(vdd), .A(_15196_), .Y(_15565_) );
NAND3X1 NAND3X1_3526 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_141_), .B(_13450_), .C(_15557_), .Y(_15566_) );
NAND2X1 NAND2X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_15381_), .B(_15561_), .Y(_15567_) );
AOI21X1 AOI21X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_15566_), .B(_15567_), .C(_15565_), .Y(_15568_) );
OAI21X1 OAI21X1_2485 ( .gnd(gnd), .vdd(vdd), .A(_15564_), .B(_15568_), .C(_15380_), .Y(_15569_) );
OAI21X1 OAI21X1_2486 ( .gnd(gnd), .vdd(vdd), .A(_15008_), .B(_15198_), .C(_15201_), .Y(_15570_) );
NAND3X1 NAND3X1_3527 ( .gnd(gnd), .vdd(vdd), .A(_15565_), .B(_15566_), .C(_15567_), .Y(_15571_) );
NAND3X1 NAND3X1_3528 ( .gnd(gnd), .vdd(vdd), .A(_15196_), .B(_15558_), .C(_15563_), .Y(_15572_) );
NAND3X1 NAND3X1_3529 ( .gnd(gnd), .vdd(vdd), .A(_15571_), .B(_15572_), .C(_15570_), .Y(_15574_) );
NAND3X1 NAND3X1_3530 ( .gnd(gnd), .vdd(vdd), .A(_15379_), .B(_15574_), .C(_15569_), .Y(_15575_) );
AOI21X1 AOI21X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_15571_), .B(_15572_), .C(_15570_), .Y(_15576_) );
NOR3X1 NOR3X1_461 ( .gnd(gnd), .vdd(vdd), .A(_15564_), .B(_15380_), .C(_15568_), .Y(_15577_) );
OAI21X1 OAI21X1_2487 ( .gnd(gnd), .vdd(vdd), .A(_15577_), .B(_15576_), .C(_16231_), .Y(_15578_) );
NAND2X1 NAND2X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_15575_), .B(_15578_), .Y(_15579_) );
NAND3X1 NAND3X1_3531 ( .gnd(gnd), .vdd(vdd), .A(_15378_), .B(_13458_), .C(_15579_), .Y(_15580_) );
OAI21X1 OAI21X1_2488 ( .gnd(gnd), .vdd(vdd), .A(_15577_), .B(_15576_), .C(_15379_), .Y(_15581_) );
NAND3X1 NAND3X1_3532 ( .gnd(gnd), .vdd(vdd), .A(_16231_), .B(_15574_), .C(_15569_), .Y(_15582_) );
NAND3X1 NAND3X1_3533 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .B(_15582_), .C(_15581_), .Y(_15583_) );
NAND2X1 NAND2X1_2003 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_157_), .B(_15583_), .Y(_15585_) );
AOI21X1 AOI21X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_15580_), .B(_15585_), .C(_15216_), .Y(_15586_) );
INVX1 INVX1_2159 ( .gnd(gnd), .vdd(vdd), .A(_15216_), .Y(_15587_) );
NAND3X1 NAND3X1_3534 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_157_), .B(_13458_), .C(_15579_), .Y(_15588_) );
NAND2X1 NAND2X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_15378_), .B(_15583_), .Y(_15589_) );
AOI21X1 AOI21X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_15588_), .B(_15589_), .C(_15587_), .Y(_15590_) );
OAI21X1 OAI21X1_2489 ( .gnd(gnd), .vdd(vdd), .A(_15586_), .B(_15590_), .C(_15377_), .Y(_15591_) );
OAI21X1 OAI21X1_2490 ( .gnd(gnd), .vdd(vdd), .A(_15218_), .B(_15006_), .C(_15223_), .Y(_15592_) );
NAND3X1 NAND3X1_3535 ( .gnd(gnd), .vdd(vdd), .A(_15587_), .B(_15588_), .C(_15589_), .Y(_15593_) );
NAND3X1 NAND3X1_3536 ( .gnd(gnd), .vdd(vdd), .A(_15216_), .B(_15580_), .C(_15585_), .Y(_15594_) );
NAND3X1 NAND3X1_3537 ( .gnd(gnd), .vdd(vdd), .A(_15593_), .B(_15594_), .C(_15592_), .Y(_15596_) );
NAND3X1 NAND3X1_3538 ( .gnd(gnd), .vdd(vdd), .A(_15376_), .B(_15596_), .C(_15591_), .Y(_15597_) );
AOI21X1 AOI21X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_15593_), .B(_15594_), .C(_15592_), .Y(_15598_) );
NOR3X1 NOR3X1_462 ( .gnd(gnd), .vdd(vdd), .A(_15586_), .B(_15377_), .C(_15590_), .Y(_15599_) );
OAI21X1 OAI21X1_2491 ( .gnd(gnd), .vdd(vdd), .A(_15599_), .B(_15598_), .C(_16315_), .Y(_15600_) );
NAND2X1 NAND2X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_15597_), .B(_15600_), .Y(_15601_) );
NAND3X1 NAND3X1_3539 ( .gnd(gnd), .vdd(vdd), .A(_15374_), .B(_13466_), .C(_15601_), .Y(_15602_) );
OAI21X1 OAI21X1_2492 ( .gnd(gnd), .vdd(vdd), .A(_15599_), .B(_15598_), .C(_15376_), .Y(_15603_) );
NAND3X1 NAND3X1_3540 ( .gnd(gnd), .vdd(vdd), .A(_16315_), .B(_15596_), .C(_15591_), .Y(_15604_) );
NAND3X1 NAND3X1_3541 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .B(_15604_), .C(_15603_), .Y(_15605_) );
NAND2X1 NAND2X1_2006 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_173_), .B(_15605_), .Y(_15607_) );
AOI21X1 AOI21X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_15602_), .B(_15607_), .C(_15229_), .Y(_15608_) );
INVX1 INVX1_2160 ( .gnd(gnd), .vdd(vdd), .A(_15229_), .Y(_15609_) );
NAND3X1 NAND3X1_3542 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_173_), .B(_13466_), .C(_15601_), .Y(_15610_) );
NAND2X1 NAND2X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_15374_), .B(_15605_), .Y(_15611_) );
AOI21X1 AOI21X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_15610_), .B(_15611_), .C(_15609_), .Y(_15612_) );
OAI21X1 OAI21X1_2493 ( .gnd(gnd), .vdd(vdd), .A(_15608_), .B(_15612_), .C(_15373_), .Y(_15613_) );
OAI21X1 OAI21X1_2494 ( .gnd(gnd), .vdd(vdd), .A(_15245_), .B(_15247_), .C(_15238_), .Y(_15614_) );
NAND3X1 NAND3X1_3543 ( .gnd(gnd), .vdd(vdd), .A(_15609_), .B(_15610_), .C(_15611_), .Y(_15615_) );
NAND3X1 NAND3X1_3544 ( .gnd(gnd), .vdd(vdd), .A(_15229_), .B(_15602_), .C(_15607_), .Y(_15616_) );
NAND3X1 NAND3X1_3545 ( .gnd(gnd), .vdd(vdd), .A(_15615_), .B(_15616_), .C(_15614_), .Y(_15618_) );
NAND3X1 NAND3X1_3546 ( .gnd(gnd), .vdd(vdd), .A(_16324_), .B(_15618_), .C(_15613_), .Y(_15619_) );
AOI21X1 AOI21X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_15615_), .B(_15616_), .C(_15614_), .Y(_15620_) );
NOR3X1 NOR3X1_463 ( .gnd(gnd), .vdd(vdd), .A(_15608_), .B(_15373_), .C(_15612_), .Y(_15621_) );
OAI21X1 OAI21X1_2495 ( .gnd(gnd), .vdd(vdd), .A(_15621_), .B(_15620_), .C(_16323_), .Y(_15622_) );
NAND2X1 NAND2X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_15619_), .B(_15622_), .Y(_15623_) );
NAND3X1 NAND3X1_3547 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_189_), .B(_13474_), .C(_15623_), .Y(_15624_) );
INVX1 INVX1_2161 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_189_), .Y(_15625_) );
OAI21X1 OAI21X1_2496 ( .gnd(gnd), .vdd(vdd), .A(_15621_), .B(_15620_), .C(_16324_), .Y(_15626_) );
NAND3X1 NAND3X1_3548 ( .gnd(gnd), .vdd(vdd), .A(_16323_), .B(_15618_), .C(_15613_), .Y(_15627_) );
NAND3X1 NAND3X1_3549 ( .gnd(gnd), .vdd(vdd), .A(_13474_), .B(_15627_), .C(_15626_), .Y(_15629_) );
NAND2X1 NAND2X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_15625_), .B(_15629_), .Y(_15630_) );
NAND3X1 NAND3X1_3550 ( .gnd(gnd), .vdd(vdd), .A(_15372_), .B(_15624_), .C(_15630_), .Y(_15631_) );
NAND3X1 NAND3X1_3551 ( .gnd(gnd), .vdd(vdd), .A(_15625_), .B(_13474_), .C(_15623_), .Y(_15632_) );
NAND2X1 NAND2X1_2010 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_189_), .B(_15629_), .Y(_15633_) );
NAND3X1 NAND3X1_3552 ( .gnd(gnd), .vdd(vdd), .A(_15254_), .B(_15632_), .C(_15633_), .Y(_15634_) );
AOI21X1 AOI21X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_15631_), .B(_15634_), .C(_15371_), .Y(_15635_) );
AOI21X1 AOI21X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_14999_), .B(_15264_), .C(_15269_), .Y(_15636_) );
AOI21X1 AOI21X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_15632_), .B(_15633_), .C(_15254_), .Y(_15637_) );
AOI21X1 AOI21X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_15624_), .B(_15630_), .C(_15372_), .Y(_15638_) );
NOR3X1 NOR3X1_464 ( .gnd(gnd), .vdd(vdd), .A(_15637_), .B(_15636_), .C(_15638_), .Y(_15640_) );
OAI21X1 OAI21X1_2497 ( .gnd(gnd), .vdd(vdd), .A(_15640_), .B(_15635_), .C(_16332_), .Y(_15641_) );
INVX1 INVX1_2162 ( .gnd(gnd), .vdd(vdd), .A(_16332_), .Y(_15642_) );
OAI21X1 OAI21X1_2498 ( .gnd(gnd), .vdd(vdd), .A(_15637_), .B(_15638_), .C(_15636_), .Y(_15643_) );
NAND3X1 NAND3X1_3553 ( .gnd(gnd), .vdd(vdd), .A(_15631_), .B(_15634_), .C(_15371_), .Y(_15644_) );
NAND3X1 NAND3X1_3554 ( .gnd(gnd), .vdd(vdd), .A(_15642_), .B(_15643_), .C(_15644_), .Y(_15645_) );
NAND2X1 NAND2X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_15645_), .B(_15641_), .Y(_15646_) );
NAND3X1 NAND3X1_3555 ( .gnd(gnd), .vdd(vdd), .A(_15370_), .B(_13482_), .C(_15646_), .Y(_15647_) );
OAI21X1 OAI21X1_2499 ( .gnd(gnd), .vdd(vdd), .A(_15640_), .B(_15635_), .C(_15642_), .Y(_15648_) );
NAND3X1 NAND3X1_3556 ( .gnd(gnd), .vdd(vdd), .A(_16332_), .B(_15643_), .C(_15644_), .Y(_15649_) );
NAND3X1 NAND3X1_3557 ( .gnd(gnd), .vdd(vdd), .A(_13482_), .B(_15649_), .C(_15648_), .Y(_15651_) );
NAND2X1 NAND2X1_2012 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_205_), .B(_15651_), .Y(_15652_) );
AOI21X1 AOI21X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_15647_), .B(_15652_), .C(_15285_), .Y(_15653_) );
INVX1 INVX1_2163 ( .gnd(gnd), .vdd(vdd), .A(_15285_), .Y(_15654_) );
NAND3X1 NAND3X1_3558 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_205_), .B(_13482_), .C(_15646_), .Y(_15655_) );
NAND2X1 NAND2X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_15370_), .B(_15651_), .Y(_15656_) );
AOI21X1 AOI21X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_15655_), .B(_15656_), .C(_15654_), .Y(_15657_) );
OAI21X1 OAI21X1_2500 ( .gnd(gnd), .vdd(vdd), .A(_15653_), .B(_15657_), .C(_15369_), .Y(_15658_) );
OAI21X1 OAI21X1_2501 ( .gnd(gnd), .vdd(vdd), .A(_15287_), .B(_14998_), .C(_15292_), .Y(_15659_) );
NAND3X1 NAND3X1_3559 ( .gnd(gnd), .vdd(vdd), .A(_15654_), .B(_15655_), .C(_15656_), .Y(_15660_) );
NAND3X1 NAND3X1_3560 ( .gnd(gnd), .vdd(vdd), .A(_15285_), .B(_15647_), .C(_15652_), .Y(_15662_) );
NAND3X1 NAND3X1_3561 ( .gnd(gnd), .vdd(vdd), .A(_15660_), .B(_15662_), .C(_15659_), .Y(_15663_) );
NAND3X1 NAND3X1_3562 ( .gnd(gnd), .vdd(vdd), .A(_16340_), .B(_15663_), .C(_15658_), .Y(_15664_) );
NAND2X1 NAND2X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_15663_), .B(_15658_), .Y(_15665_) );
AOI21X1 AOI21X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_16341_), .B(_15665_), .C(_13491_), .Y(_15666_) );
NAND3X1 NAND3X1_3563 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_221_), .B(_15664_), .C(_15666_), .Y(_15667_) );
INVX1 INVX1_2164 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_221_), .Y(_15668_) );
AOI21X1 AOI21X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_15660_), .B(_15662_), .C(_15659_), .Y(_15669_) );
NOR3X1 NOR3X1_465 ( .gnd(gnd), .vdd(vdd), .A(_15369_), .B(_15653_), .C(_15657_), .Y(_15670_) );
OAI21X1 OAI21X1_2502 ( .gnd(gnd), .vdd(vdd), .A(_15670_), .B(_15669_), .C(_16341_), .Y(_15671_) );
NAND3X1 NAND3X1_3564 ( .gnd(gnd), .vdd(vdd), .A(_13490_), .B(_15664_), .C(_15671_), .Y(_15673_) );
NAND2X1 NAND2X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_15668_), .B(_15673_), .Y(_15674_) );
NAND3X1 NAND3X1_3565 ( .gnd(gnd), .vdd(vdd), .A(_15368_), .B(_15667_), .C(_15674_), .Y(_15675_) );
NAND3X1 NAND3X1_3566 ( .gnd(gnd), .vdd(vdd), .A(_15668_), .B(_15664_), .C(_15666_), .Y(_15676_) );
NAND2X1 NAND2X1_2016 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_221_), .B(_15673_), .Y(_15677_) );
NAND3X1 NAND3X1_3567 ( .gnd(gnd), .vdd(vdd), .A(_15308_), .B(_15676_), .C(_15677_), .Y(_15678_) );
AOI21X1 AOI21X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_15675_), .B(_15678_), .C(_15367_), .Y(_15679_) );
AOI21X1 AOI21X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_15315_), .B(_15317_), .C(_15307_), .Y(_15680_) );
AOI21X1 AOI21X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_15676_), .B(_15677_), .C(_15308_), .Y(_15681_) );
AOI21X1 AOI21X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_15667_), .B(_15674_), .C(_15368_), .Y(_15682_) );
NOR3X1 NOR3X1_466 ( .gnd(gnd), .vdd(vdd), .A(_15681_), .B(_15680_), .C(_15682_), .Y(_15684_) );
OAI21X1 OAI21X1_2503 ( .gnd(gnd), .vdd(vdd), .A(_15684_), .B(_15679_), .C(_16349_), .Y(_15685_) );
INVX1 INVX1_2165 ( .gnd(gnd), .vdd(vdd), .A(_16349_), .Y(_15686_) );
OAI21X1 OAI21X1_2504 ( .gnd(gnd), .vdd(vdd), .A(_15681_), .B(_15682_), .C(_15680_), .Y(_15687_) );
NAND3X1 NAND3X1_3568 ( .gnd(gnd), .vdd(vdd), .A(_15675_), .B(_15678_), .C(_15367_), .Y(_15688_) );
NAND3X1 NAND3X1_3569 ( .gnd(gnd), .vdd(vdd), .A(_15686_), .B(_15688_), .C(_15687_), .Y(_15689_) );
NAND2X1 NAND2X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_15689_), .B(_15685_), .Y(_15690_) );
NAND3X1 NAND3X1_3570 ( .gnd(gnd), .vdd(vdd), .A(_15366_), .B(_13498_), .C(_15690_), .Y(_15691_) );
OAI21X1 OAI21X1_2505 ( .gnd(gnd), .vdd(vdd), .A(_15684_), .B(_15679_), .C(_15686_), .Y(_15692_) );
NAND3X1 NAND3X1_3571 ( .gnd(gnd), .vdd(vdd), .A(_16349_), .B(_15688_), .C(_15687_), .Y(_15693_) );
NAND3X1 NAND3X1_3572 ( .gnd(gnd), .vdd(vdd), .A(_13498_), .B(_15693_), .C(_15692_), .Y(_15695_) );
NAND2X1 NAND2X1_2018 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_237_), .B(_15695_), .Y(_15696_) );
AOI21X1 AOI21X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_15691_), .B(_15696_), .C(_15323_), .Y(_15697_) );
INVX1 INVX1_2166 ( .gnd(gnd), .vdd(vdd), .A(_15323_), .Y(_15698_) );
NAND3X1 NAND3X1_3573 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_237_), .B(_13498_), .C(_15690_), .Y(_15699_) );
NAND2X1 NAND2X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_15366_), .B(_15695_), .Y(_15700_) );
AOI21X1 AOI21X1_2220 ( .gnd(gnd), .vdd(vdd), .A(_15699_), .B(_15700_), .C(_15698_), .Y(_15701_) );
OAI21X1 OAI21X1_2506 ( .gnd(gnd), .vdd(vdd), .A(_15697_), .B(_15701_), .C(_15365_), .Y(_15702_) );
OAI21X1 OAI21X1_2507 ( .gnd(gnd), .vdd(vdd), .A(_15338_), .B(_15345_), .C(_15331_), .Y(_15703_) );
NAND3X1 NAND3X1_3574 ( .gnd(gnd), .vdd(vdd), .A(_15698_), .B(_15699_), .C(_15700_), .Y(_15704_) );
NAND3X1 NAND3X1_3575 ( .gnd(gnd), .vdd(vdd), .A(_15323_), .B(_15691_), .C(_15696_), .Y(_15706_) );
NAND3X1 NAND3X1_3576 ( .gnd(gnd), .vdd(vdd), .A(_15704_), .B(_15706_), .C(_15703_), .Y(_15707_) );
NAND3X1 NAND3X1_3577 ( .gnd(gnd), .vdd(vdd), .A(_16546_), .B(_15702_), .C(_15707_), .Y(_15708_) );
AOI21X1 AOI21X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_15704_), .B(_15706_), .C(_15703_), .Y(_15709_) );
NOR3X1 NOR3X1_467 ( .gnd(gnd), .vdd(vdd), .A(_15697_), .B(_15365_), .C(_15701_), .Y(_15710_) );
OAI21X1 OAI21X1_2508 ( .gnd(gnd), .vdd(vdd), .A(_15710_), .B(_15709_), .C(_16357_), .Y(_15711_) );
NAND2X1 NAND2X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_15708_), .B(_15711_), .Y(_15712_) );
NAND3X1 NAND3X1_3578 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_253_), .B(_13506_), .C(_15712_), .Y(_15713_) );
INVX1 INVX1_2167 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_253_), .Y(_15714_) );
OAI21X1 OAI21X1_2509 ( .gnd(gnd), .vdd(vdd), .A(_15710_), .B(_15709_), .C(_16546_), .Y(_15715_) );
NAND3X1 NAND3X1_3579 ( .gnd(gnd), .vdd(vdd), .A(_16357_), .B(_15702_), .C(_15707_), .Y(_15717_) );
NAND3X1 NAND3X1_3580 ( .gnd(gnd), .vdd(vdd), .A(_13506_), .B(_15717_), .C(_15715_), .Y(_15718_) );
NAND2X1 NAND2X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_15714_), .B(_15718_), .Y(_15719_) );
NAND3X1 NAND3X1_3581 ( .gnd(gnd), .vdd(vdd), .A(_15363_), .B(_15713_), .C(_15719_), .Y(_15720_) );
INVX1 INVX1_2168 ( .gnd(gnd), .vdd(vdd), .A(_15363_), .Y(_15721_) );
NAND2X1 NAND2X1_2022 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_253_), .B(_15718_), .Y(_15722_) );
OR2X2 OR2X2_363 ( .gnd(gnd), .vdd(vdd), .A(_15718_), .B(module_3_W_253_), .Y(_15723_) );
NAND3X1 NAND3X1_3582 ( .gnd(gnd), .vdd(vdd), .A(_15721_), .B(_15722_), .C(_15723_), .Y(_15724_) );
NAND2X1 NAND2X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_15720_), .B(_15724_), .Y(_15725_) );
XNOR2X1 XNOR2X1_402 ( .gnd(gnd), .vdd(vdd), .A(_15725_), .B(_15361_), .Y(module_3_H_21_) );
AOI21X1 AOI21X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_15713_), .B(_15719_), .C(_15363_), .Y(_15727_) );
AOI21X1 AOI21X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_15361_), .B(_15720_), .C(_15727_), .Y(_15728_) );
INVX1 INVX1_2169 ( .gnd(gnd), .vdd(vdd), .A(_15728_), .Y(_15729_) );
INVX1 INVX1_2170 ( .gnd(gnd), .vdd(vdd), .A(_15722_), .Y(_15730_) );
OAI21X1 OAI21X1_2510 ( .gnd(gnd), .vdd(vdd), .A(_15701_), .B(_15365_), .C(_15704_), .Y(_15731_) );
OAI21X1 OAI21X1_2511 ( .gnd(gnd), .vdd(vdd), .A(_15682_), .B(_15680_), .C(_15675_), .Y(_15732_) );
OAI21X1 OAI21X1_2512 ( .gnd(gnd), .vdd(vdd), .A(_15369_), .B(_15657_), .C(_15660_), .Y(_15733_) );
OAI21X1 OAI21X1_2513 ( .gnd(gnd), .vdd(vdd), .A(_15638_), .B(_15636_), .C(_15631_), .Y(_15734_) );
INVX1 INVX1_2171 ( .gnd(gnd), .vdd(vdd), .A(_15734_), .Y(_15735_) );
INVX1 INVX1_2172 ( .gnd(gnd), .vdd(vdd), .A(_15632_), .Y(_15736_) );
OAI21X1 OAI21X1_2514 ( .gnd(gnd), .vdd(vdd), .A(_15612_), .B(_15373_), .C(_15615_), .Y(_15738_) );
INVX1 INVX1_2173 ( .gnd(gnd), .vdd(vdd), .A(_15738_), .Y(_15739_) );
INVX1 INVX1_2174 ( .gnd(gnd), .vdd(vdd), .A(_15602_), .Y(_15740_) );
OAI21X1 OAI21X1_2515 ( .gnd(gnd), .vdd(vdd), .A(_15590_), .B(_15377_), .C(_15593_), .Y(_15741_) );
INVX1 INVX1_2175 ( .gnd(gnd), .vdd(vdd), .A(_15741_), .Y(_15742_) );
INVX1 INVX1_2176 ( .gnd(gnd), .vdd(vdd), .A(_15580_), .Y(_15743_) );
OAI21X1 OAI21X1_2516 ( .gnd(gnd), .vdd(vdd), .A(_15568_), .B(_15380_), .C(_15571_), .Y(_15744_) );
NAND2X1 NAND2X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_15542_), .B(_15555_), .Y(_15745_) );
INVX1 INVX1_2177 ( .gnd(gnd), .vdd(vdd), .A(_15745_), .Y(_15746_) );
NAND2X1 NAND2X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_15527_), .B(_15530_), .Y(_15747_) );
NAND2X1 NAND2X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_15506_), .B(_15509_), .Y(_15749_) );
NAND2X1 NAND2X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_15486_), .B(_15488_), .Y(_15750_) );
NAND2X1 NAND2X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_15457_), .B(_15471_), .Y(_15751_) );
NAND2X1 NAND2X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_15443_), .B(_15445_), .Y(_15752_) );
OAI21X1 OAI21X1_2517 ( .gnd(gnd), .vdd(vdd), .A(_15421_), .B(_15422_), .C(_15418_), .Y(_15753_) );
INVX1 INVX1_2178 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_30_), .Y(_15754_) );
NOR2X1 NOR2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_12_), .B(module_3_W_13_), .Y(_15755_) );
XNOR2X1 XNOR2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_15755_), .B(module_3_W_14_), .Y(_15756_) );
XNOR2X1 XNOR2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_13896_), .B(module_3_W_10_), .Y(_15757_) );
XNOR2X1 XNOR2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_15757_), .B(_15756_), .Y(_15758_) );
OR2X2 OR2X2_364 ( .gnd(gnd), .vdd(vdd), .A(_15758_), .B(_15754_), .Y(_15760_) );
NAND2X1 NAND2X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_15754_), .B(_15758_), .Y(_15761_) );
NAND2X1 NAND2X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_15761_), .B(_15760_), .Y(_15762_) );
XNOR2X1 XNOR2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_15762_), .B(_15414_), .Y(_15763_) );
XOR2X1 XOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_15763_), .B(_15753_), .Y(_15764_) );
XNOR2X1 XNOR2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_13920_), .B(_13955_), .Y(_15765_) );
XOR2X1 XOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_15764_), .B(_15765_), .Y(_15766_) );
NAND2X1 NAND2X1_2032 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf3_), .B(_15766_), .Y(_15767_) );
INVX1 INVX1_2179 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf2_), .Y(_15768_) );
XNOR2X1 XNOR2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_15764_), .B(_15765_), .Y(_15769_) );
NAND2X1 NAND2X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_15768_), .B(_15769_), .Y(_15771_) );
NAND3X1 NAND3X1_3583 ( .gnd(gnd), .vdd(vdd), .A(_15438_), .B(_15771_), .C(_15767_), .Y(_15772_) );
NAND2X1 NAND2X1_2034 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf1_), .B(_15769_), .Y(_15773_) );
NAND2X1 NAND2X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_15768_), .B(_15766_), .Y(_15774_) );
NAND3X1 NAND3X1_3584 ( .gnd(gnd), .vdd(vdd), .A(_15435_), .B(_15773_), .C(_15774_), .Y(_15775_) );
NAND3X1 NAND3X1_3585 ( .gnd(gnd), .vdd(vdd), .A(_15752_), .B(_15772_), .C(_15775_), .Y(_15776_) );
AOI21X1 AOI21X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_15772_), .B(_15775_), .C(_15752_), .Y(_15777_) );
INVX1 INVX1_2180 ( .gnd(gnd), .vdd(vdd), .A(_15777_), .Y(_15778_) );
XNOR2X1 XNOR2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_13990_), .B(_13941_), .Y(_15779_) );
NAND3X1 NAND3X1_3586 ( .gnd(gnd), .vdd(vdd), .A(_15776_), .B(_15779_), .C(_15778_), .Y(_15780_) );
INVX1 INVX1_2181 ( .gnd(gnd), .vdd(vdd), .A(_15776_), .Y(_15782_) );
INVX1 INVX1_2182 ( .gnd(gnd), .vdd(vdd), .A(_15779_), .Y(_15783_) );
OAI21X1 OAI21X1_2518 ( .gnd(gnd), .vdd(vdd), .A(_15782_), .B(_15777_), .C(_15783_), .Y(_15784_) );
NAND3X1 NAND3X1_3587 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf0_), .B(_15780_), .C(_15784_), .Y(_15785_) );
INVX1 INVX1_2183 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf3_), .Y(_15786_) );
OAI21X1 OAI21X1_2519 ( .gnd(gnd), .vdd(vdd), .A(_15782_), .B(_15777_), .C(_15779_), .Y(_15787_) );
NAND3X1 NAND3X1_3588 ( .gnd(gnd), .vdd(vdd), .A(_15776_), .B(_15783_), .C(_15778_), .Y(_15788_) );
NAND3X1 NAND3X1_3589 ( .gnd(gnd), .vdd(vdd), .A(_15786_), .B(_15788_), .C(_15787_), .Y(_15789_) );
NAND3X1 NAND3X1_3590 ( .gnd(gnd), .vdd(vdd), .A(_15460_), .B(_15785_), .C(_15789_), .Y(_15790_) );
NAND3X1 NAND3X1_3591 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf2_), .B(_15788_), .C(_15787_), .Y(_15791_) );
NAND3X1 NAND3X1_3592 ( .gnd(gnd), .vdd(vdd), .A(_15786_), .B(_15780_), .C(_15784_), .Y(_15793_) );
NAND3X1 NAND3X1_3593 ( .gnd(gnd), .vdd(vdd), .A(_15456_), .B(_15791_), .C(_15793_), .Y(_15794_) );
NAND3X1 NAND3X1_3594 ( .gnd(gnd), .vdd(vdd), .A(_15751_), .B(_15790_), .C(_15794_), .Y(_15795_) );
INVX1 INVX1_2184 ( .gnd(gnd), .vdd(vdd), .A(_15751_), .Y(_15796_) );
NAND3X1 NAND3X1_3595 ( .gnd(gnd), .vdd(vdd), .A(_15460_), .B(_15791_), .C(_15793_), .Y(_15797_) );
NAND3X1 NAND3X1_3596 ( .gnd(gnd), .vdd(vdd), .A(_15456_), .B(_15785_), .C(_15789_), .Y(_15798_) );
NAND3X1 NAND3X1_3597 ( .gnd(gnd), .vdd(vdd), .A(_15796_), .B(_15797_), .C(_15798_), .Y(_15799_) );
XNOR2X1 XNOR2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_14028_), .B(_13978_), .Y(_15800_) );
NAND3X1 NAND3X1_3598 ( .gnd(gnd), .vdd(vdd), .A(_15800_), .B(_15795_), .C(_15799_), .Y(_15801_) );
AOI21X1 AOI21X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_15797_), .B(_15798_), .C(_15796_), .Y(_15802_) );
AOI21X1 AOI21X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_15790_), .B(_15794_), .C(_15751_), .Y(_15804_) );
INVX1 INVX1_2185 ( .gnd(gnd), .vdd(vdd), .A(_15800_), .Y(_15805_) );
OAI21X1 OAI21X1_2520 ( .gnd(gnd), .vdd(vdd), .A(_15802_), .B(_15804_), .C(_15805_), .Y(_15806_) );
NAND3X1 NAND3X1_3599 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf1_), .B(_15801_), .C(_15806_), .Y(_15807_) );
INVX1 INVX1_2186 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf0_), .Y(_15808_) );
OAI21X1 OAI21X1_2521 ( .gnd(gnd), .vdd(vdd), .A(_15802_), .B(_15804_), .C(_15800_), .Y(_15809_) );
NAND3X1 NAND3X1_3600 ( .gnd(gnd), .vdd(vdd), .A(_15805_), .B(_15795_), .C(_15799_), .Y(_15810_) );
NAND3X1 NAND3X1_3601 ( .gnd(gnd), .vdd(vdd), .A(_15808_), .B(_15810_), .C(_15809_), .Y(_15811_) );
NAND3X1 NAND3X1_3602 ( .gnd(gnd), .vdd(vdd), .A(_15481_), .B(_15807_), .C(_15811_), .Y(_15812_) );
NAND3X1 NAND3X1_3603 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf4_), .B(_15810_), .C(_15809_), .Y(_15813_) );
NAND3X1 NAND3X1_3604 ( .gnd(gnd), .vdd(vdd), .A(_15808_), .B(_15801_), .C(_15806_), .Y(_15815_) );
NAND3X1 NAND3X1_3605 ( .gnd(gnd), .vdd(vdd), .A(_15478_), .B(_15813_), .C(_15815_), .Y(_15816_) );
NAND3X1 NAND3X1_3606 ( .gnd(gnd), .vdd(vdd), .A(_15750_), .B(_15812_), .C(_15816_), .Y(_15817_) );
INVX1 INVX1_2187 ( .gnd(gnd), .vdd(vdd), .A(_15750_), .Y(_15818_) );
NAND3X1 NAND3X1_3607 ( .gnd(gnd), .vdd(vdd), .A(_15481_), .B(_15813_), .C(_15815_), .Y(_15819_) );
NAND3X1 NAND3X1_3608 ( .gnd(gnd), .vdd(vdd), .A(_15478_), .B(_15807_), .C(_15811_), .Y(_15820_) );
NAND3X1 NAND3X1_3609 ( .gnd(gnd), .vdd(vdd), .A(_15818_), .B(_15819_), .C(_15820_), .Y(_15821_) );
XNOR2X1 XNOR2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_14067_), .B(_16644_), .Y(_15822_) );
NAND3X1 NAND3X1_3610 ( .gnd(gnd), .vdd(vdd), .A(_15822_), .B(_15817_), .C(_15821_), .Y(_15823_) );
AOI21X1 AOI21X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_15819_), .B(_15820_), .C(_15818_), .Y(_15824_) );
AOI21X1 AOI21X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_15812_), .B(_15816_), .C(_15750_), .Y(_15826_) );
INVX1 INVX1_2188 ( .gnd(gnd), .vdd(vdd), .A(_15822_), .Y(_15827_) );
OAI21X1 OAI21X1_2522 ( .gnd(gnd), .vdd(vdd), .A(_15824_), .B(_15826_), .C(_15827_), .Y(_15828_) );
NAND3X1 NAND3X1_3611 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf0_), .B(_15823_), .C(_15828_), .Y(_15829_) );
INVX1 INVX1_2189 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf3_), .Y(_15830_) );
OAI21X1 OAI21X1_2523 ( .gnd(gnd), .vdd(vdd), .A(_15824_), .B(_15826_), .C(_15822_), .Y(_15831_) );
NAND3X1 NAND3X1_3612 ( .gnd(gnd), .vdd(vdd), .A(_15827_), .B(_15817_), .C(_15821_), .Y(_15832_) );
NAND3X1 NAND3X1_3613 ( .gnd(gnd), .vdd(vdd), .A(_15830_), .B(_15832_), .C(_15831_), .Y(_15833_) );
NAND3X1 NAND3X1_3614 ( .gnd(gnd), .vdd(vdd), .A(_15502_), .B(_15829_), .C(_15833_), .Y(_15834_) );
NAND3X1 NAND3X1_3615 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf2_), .B(_15832_), .C(_15831_), .Y(_15835_) );
NAND3X1 NAND3X1_3616 ( .gnd(gnd), .vdd(vdd), .A(_15830_), .B(_15823_), .C(_15828_), .Y(_15837_) );
NAND3X1 NAND3X1_3617 ( .gnd(gnd), .vdd(vdd), .A(_15499_), .B(_15835_), .C(_15837_), .Y(_15838_) );
NAND3X1 NAND3X1_3618 ( .gnd(gnd), .vdd(vdd), .A(_15749_), .B(_15834_), .C(_15838_), .Y(_15839_) );
INVX2 INVX2_535 ( .gnd(gnd), .vdd(vdd), .A(_15749_), .Y(_15840_) );
AOI21X1 AOI21X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_15835_), .B(_15837_), .C(_15499_), .Y(_15841_) );
AOI21X1 AOI21X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_15829_), .B(_15833_), .C(_15502_), .Y(_15842_) );
OAI21X1 OAI21X1_2524 ( .gnd(gnd), .vdd(vdd), .A(_15841_), .B(_15842_), .C(_15840_), .Y(_15843_) );
XOR2X1 XOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_14108_), .B(_14069_), .Y(_15844_) );
NAND3X1 NAND3X1_3619 ( .gnd(gnd), .vdd(vdd), .A(_15839_), .B(_15844_), .C(_15843_), .Y(_15845_) );
NOR3X1 NOR3X1_468 ( .gnd(gnd), .vdd(vdd), .A(_15841_), .B(_15840_), .C(_15842_), .Y(_15846_) );
AOI21X1 AOI21X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_15834_), .B(_15838_), .C(_15749_), .Y(_15848_) );
INVX1 INVX1_2190 ( .gnd(gnd), .vdd(vdd), .A(_15844_), .Y(_15849_) );
OAI21X1 OAI21X1_2525 ( .gnd(gnd), .vdd(vdd), .A(_15846_), .B(_15848_), .C(_15849_), .Y(_15850_) );
NAND3X1 NAND3X1_3620 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf1_), .B(_15845_), .C(_15850_), .Y(_15851_) );
INVX1 INVX1_2191 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf0_), .Y(_15852_) );
OAI21X1 OAI21X1_2526 ( .gnd(gnd), .vdd(vdd), .A(_15846_), .B(_15848_), .C(_15844_), .Y(_15853_) );
NAND3X1 NAND3X1_3621 ( .gnd(gnd), .vdd(vdd), .A(_15839_), .B(_15849_), .C(_15843_), .Y(_15854_) );
NAND3X1 NAND3X1_3622 ( .gnd(gnd), .vdd(vdd), .A(_15852_), .B(_15854_), .C(_15853_), .Y(_15855_) );
NAND3X1 NAND3X1_3623 ( .gnd(gnd), .vdd(vdd), .A(_15523_), .B(_15851_), .C(_15855_), .Y(_15856_) );
NAND3X1 NAND3X1_3624 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf4_), .B(_15854_), .C(_15853_), .Y(_15857_) );
NAND3X1 NAND3X1_3625 ( .gnd(gnd), .vdd(vdd), .A(_15852_), .B(_15845_), .C(_15850_), .Y(_15859_) );
NAND3X1 NAND3X1_3626 ( .gnd(gnd), .vdd(vdd), .A(_15520_), .B(_15857_), .C(_15859_), .Y(_15860_) );
NAND3X1 NAND3X1_3627 ( .gnd(gnd), .vdd(vdd), .A(_15747_), .B(_15856_), .C(_15860_), .Y(_15861_) );
INVX1 INVX1_2192 ( .gnd(gnd), .vdd(vdd), .A(_15747_), .Y(_15862_) );
NAND3X1 NAND3X1_3628 ( .gnd(gnd), .vdd(vdd), .A(_15523_), .B(_15857_), .C(_15859_), .Y(_15863_) );
NAND3X1 NAND3X1_3629 ( .gnd(gnd), .vdd(vdd), .A(_15520_), .B(_15851_), .C(_15855_), .Y(_15864_) );
NAND3X1 NAND3X1_3630 ( .gnd(gnd), .vdd(vdd), .A(_15862_), .B(_15863_), .C(_15864_), .Y(_15865_) );
XOR2X1 XOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_14148_), .B(_14110_), .Y(_15866_) );
INVX1 INVX1_2193 ( .gnd(gnd), .vdd(vdd), .A(_15866_), .Y(_15867_) );
NAND3X1 NAND3X1_3631 ( .gnd(gnd), .vdd(vdd), .A(_15867_), .B(_15861_), .C(_15865_), .Y(_15868_) );
AOI21X1 AOI21X1_2232 ( .gnd(gnd), .vdd(vdd), .A(_15863_), .B(_15864_), .C(_15862_), .Y(_15870_) );
AOI21X1 AOI21X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_15856_), .B(_15860_), .C(_15747_), .Y(_15871_) );
OAI21X1 OAI21X1_2527 ( .gnd(gnd), .vdd(vdd), .A(_15870_), .B(_15871_), .C(_15866_), .Y(_15872_) );
NAND3X1 NAND3X1_3632 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf3_), .B(_15868_), .C(_15872_), .Y(_15873_) );
INVX1 INVX1_2194 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf2_), .Y(_15874_) );
NAND3X1 NAND3X1_3633 ( .gnd(gnd), .vdd(vdd), .A(_15866_), .B(_15861_), .C(_15865_), .Y(_15875_) );
OAI21X1 OAI21X1_2528 ( .gnd(gnd), .vdd(vdd), .A(_15870_), .B(_15871_), .C(_15867_), .Y(_15876_) );
NAND3X1 NAND3X1_3634 ( .gnd(gnd), .vdd(vdd), .A(_15874_), .B(_15875_), .C(_15876_), .Y(_15877_) );
NAND3X1 NAND3X1_3635 ( .gnd(gnd), .vdd(vdd), .A(_15545_), .B(_15873_), .C(_15877_), .Y(_15878_) );
NAND3X1 NAND3X1_3636 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf1_), .B(_15875_), .C(_15876_), .Y(_15879_) );
NAND3X1 NAND3X1_3637 ( .gnd(gnd), .vdd(vdd), .A(_15874_), .B(_15868_), .C(_15872_), .Y(_15881_) );
NAND3X1 NAND3X1_3638 ( .gnd(gnd), .vdd(vdd), .A(_15541_), .B(_15879_), .C(_15881_), .Y(_15882_) );
AOI21X1 AOI21X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_15878_), .B(_15882_), .C(_15746_), .Y(_15883_) );
NAND3X1 NAND3X1_3639 ( .gnd(gnd), .vdd(vdd), .A(_15545_), .B(_15879_), .C(_15881_), .Y(_15884_) );
NAND3X1 NAND3X1_3640 ( .gnd(gnd), .vdd(vdd), .A(_15541_), .B(_15873_), .C(_15877_), .Y(_15885_) );
AOI21X1 AOI21X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_15884_), .B(_15885_), .C(_15745_), .Y(_15886_) );
OAI21X1 OAI21X1_2529 ( .gnd(gnd), .vdd(vdd), .A(_15883_), .B(_15886_), .C(_14150_), .Y(_15887_) );
INVX1 INVX1_2195 ( .gnd(gnd), .vdd(vdd), .A(_14150_), .Y(_15888_) );
NAND3X1 NAND3X1_3641 ( .gnd(gnd), .vdd(vdd), .A(_15745_), .B(_15884_), .C(_15885_), .Y(_15889_) );
NAND3X1 NAND3X1_3642 ( .gnd(gnd), .vdd(vdd), .A(_15878_), .B(_15882_), .C(_15746_), .Y(_15890_) );
NAND3X1 NAND3X1_3643 ( .gnd(gnd), .vdd(vdd), .A(_15888_), .B(_15889_), .C(_15890_), .Y(_15892_) );
NAND3X1 NAND3X1_3644 ( .gnd(gnd), .vdd(vdd), .A(_14189_), .B(_15892_), .C(_15887_), .Y(_15893_) );
NAND2X1 NAND2X1_2036 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_142_), .B(_15893_), .Y(_15894_) );
INVX1 INVX1_2196 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_142_), .Y(_15895_) );
OAI21X1 OAI21X1_2530 ( .gnd(gnd), .vdd(vdd), .A(_15883_), .B(_15886_), .C(_15888_), .Y(_15896_) );
NAND3X1 NAND3X1_3645 ( .gnd(gnd), .vdd(vdd), .A(_14150_), .B(_15889_), .C(_15890_), .Y(_15897_) );
NAND2X1 NAND2X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_15897_), .B(_15896_), .Y(_15898_) );
NAND3X1 NAND3X1_3646 ( .gnd(gnd), .vdd(vdd), .A(_15895_), .B(_14189_), .C(_15898_), .Y(_15899_) );
NAND3X1 NAND3X1_3647 ( .gnd(gnd), .vdd(vdd), .A(_15558_), .B(_15899_), .C(_15894_), .Y(_15900_) );
INVX1 INVX1_2197 ( .gnd(gnd), .vdd(vdd), .A(_15558_), .Y(_15901_) );
NAND3X1 NAND3X1_3648 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_142_), .B(_14189_), .C(_15898_), .Y(_15903_) );
NAND2X1 NAND2X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_15895_), .B(_15893_), .Y(_15904_) );
NAND3X1 NAND3X1_3649 ( .gnd(gnd), .vdd(vdd), .A(_15901_), .B(_15903_), .C(_15904_), .Y(_15905_) );
NAND3X1 NAND3X1_3650 ( .gnd(gnd), .vdd(vdd), .A(_15744_), .B(_15900_), .C(_15905_), .Y(_15906_) );
INVX1 INVX1_2198 ( .gnd(gnd), .vdd(vdd), .A(_15744_), .Y(_15907_) );
NAND3X1 NAND3X1_3651 ( .gnd(gnd), .vdd(vdd), .A(_15901_), .B(_15899_), .C(_15894_), .Y(_15908_) );
NAND3X1 NAND3X1_3652 ( .gnd(gnd), .vdd(vdd), .A(_15558_), .B(_15903_), .C(_15904_), .Y(_15909_) );
NAND3X1 NAND3X1_3653 ( .gnd(gnd), .vdd(vdd), .A(_15907_), .B(_15908_), .C(_15909_), .Y(_15910_) );
NAND3X1 NAND3X1_3654 ( .gnd(gnd), .vdd(vdd), .A(_13877_), .B(_15906_), .C(_15910_), .Y(_15911_) );
AOI21X1 AOI21X1_2236 ( .gnd(gnd), .vdd(vdd), .A(_15908_), .B(_15909_), .C(_15907_), .Y(_15912_) );
AOI21X1 AOI21X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .B(_15905_), .C(_15744_), .Y(_15914_) );
OAI21X1 OAI21X1_2531 ( .gnd(gnd), .vdd(vdd), .A(_15912_), .B(_15914_), .C(_13876_), .Y(_15915_) );
NAND3X1 NAND3X1_3655 ( .gnd(gnd), .vdd(vdd), .A(_14223_), .B(_15911_), .C(_15915_), .Y(_15916_) );
NAND2X1 NAND2X1_2039 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_158_), .B(_15916_), .Y(_15917_) );
INVX1 INVX1_2199 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_158_), .Y(_15918_) );
NAND2X1 NAND2X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_15906_), .B(_15910_), .Y(_15919_) );
AOI21X1 AOI21X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_13876_), .B(_15919_), .C(_14224_), .Y(_15920_) );
NAND3X1 NAND3X1_3656 ( .gnd(gnd), .vdd(vdd), .A(_15918_), .B(_15911_), .C(_15920_), .Y(_15921_) );
NAND3X1 NAND3X1_3657 ( .gnd(gnd), .vdd(vdd), .A(_15743_), .B(_15921_), .C(_15917_), .Y(_15922_) );
NAND3X1 NAND3X1_3658 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_158_), .B(_15911_), .C(_15920_), .Y(_15923_) );
NAND2X1 NAND2X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_15918_), .B(_15916_), .Y(_15925_) );
NAND3X1 NAND3X1_3659 ( .gnd(gnd), .vdd(vdd), .A(_15580_), .B(_15923_), .C(_15925_), .Y(_15926_) );
AOI21X1 AOI21X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_15922_), .B(_15926_), .C(_15742_), .Y(_15927_) );
NAND3X1 NAND3X1_3660 ( .gnd(gnd), .vdd(vdd), .A(_15580_), .B(_15921_), .C(_15917_), .Y(_15928_) );
NAND3X1 NAND3X1_3661 ( .gnd(gnd), .vdd(vdd), .A(_15743_), .B(_15923_), .C(_15925_), .Y(_15929_) );
AOI21X1 AOI21X1_2240 ( .gnd(gnd), .vdd(vdd), .A(_15928_), .B(_15929_), .C(_15741_), .Y(_15930_) );
OAI21X1 OAI21X1_2532 ( .gnd(gnd), .vdd(vdd), .A(_15927_), .B(_15930_), .C(_16489_), .Y(_15931_) );
NAND3X1 NAND3X1_3662 ( .gnd(gnd), .vdd(vdd), .A(_15741_), .B(_15928_), .C(_15929_), .Y(_15932_) );
NAND3X1 NAND3X1_3663 ( .gnd(gnd), .vdd(vdd), .A(_15742_), .B(_15922_), .C(_15926_), .Y(_15933_) );
NAND3X1 NAND3X1_3664 ( .gnd(gnd), .vdd(vdd), .A(_16702_), .B(_15932_), .C(_15933_), .Y(_15934_) );
NAND3X1 NAND3X1_3665 ( .gnd(gnd), .vdd(vdd), .A(_14258_), .B(_15934_), .C(_15931_), .Y(_15936_) );
NAND2X1 NAND2X1_2042 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_174_), .B(_15936_), .Y(_15937_) );
INVX1 INVX1_2200 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_174_), .Y(_15938_) );
OAI21X1 OAI21X1_2533 ( .gnd(gnd), .vdd(vdd), .A(_15927_), .B(_15930_), .C(_16702_), .Y(_15939_) );
NAND3X1 NAND3X1_3666 ( .gnd(gnd), .vdd(vdd), .A(_16489_), .B(_15932_), .C(_15933_), .Y(_15940_) );
NAND2X1 NAND2X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_15940_), .B(_15939_), .Y(_15941_) );
NAND3X1 NAND3X1_3667 ( .gnd(gnd), .vdd(vdd), .A(_15938_), .B(_14258_), .C(_15941_), .Y(_15942_) );
NAND3X1 NAND3X1_3668 ( .gnd(gnd), .vdd(vdd), .A(_15740_), .B(_15942_), .C(_15937_), .Y(_15943_) );
NAND3X1 NAND3X1_3669 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_174_), .B(_14258_), .C(_15941_), .Y(_15944_) );
NAND2X1 NAND2X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_15938_), .B(_15936_), .Y(_15945_) );
NAND3X1 NAND3X1_3670 ( .gnd(gnd), .vdd(vdd), .A(_15602_), .B(_15944_), .C(_15945_), .Y(_15947_) );
AOI21X1 AOI21X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_15943_), .B(_15947_), .C(_15739_), .Y(_15948_) );
NAND3X1 NAND3X1_3671 ( .gnd(gnd), .vdd(vdd), .A(_15602_), .B(_15942_), .C(_15937_), .Y(_15949_) );
NAND3X1 NAND3X1_3672 ( .gnd(gnd), .vdd(vdd), .A(_15740_), .B(_15944_), .C(_15945_), .Y(_15950_) );
AOI21X1 AOI21X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_15949_), .B(_15950_), .C(_15738_), .Y(_15951_) );
OAI21X1 OAI21X1_2534 ( .gnd(gnd), .vdd(vdd), .A(_15951_), .B(_15948_), .C(_16499_), .Y(_15952_) );
NAND3X1 NAND3X1_3673 ( .gnd(gnd), .vdd(vdd), .A(_15738_), .B(_15949_), .C(_15950_), .Y(_15953_) );
NAND3X1 NAND3X1_3674 ( .gnd(gnd), .vdd(vdd), .A(_15943_), .B(_15739_), .C(_15947_), .Y(_15954_) );
NAND3X1 NAND3X1_3675 ( .gnd(gnd), .vdd(vdd), .A(_13871_), .B(_15953_), .C(_15954_), .Y(_15955_) );
NAND3X1 NAND3X1_3676 ( .gnd(gnd), .vdd(vdd), .A(_14296_), .B(_15955_), .C(_15952_), .Y(_15956_) );
NAND2X1 NAND2X1_2045 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_190_), .B(_15956_), .Y(_15958_) );
INVX1 INVX1_2201 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_190_), .Y(_15959_) );
OAI21X1 OAI21X1_2535 ( .gnd(gnd), .vdd(vdd), .A(_15951_), .B(_15948_), .C(_13871_), .Y(_15960_) );
NAND3X1 NAND3X1_3677 ( .gnd(gnd), .vdd(vdd), .A(_16499_), .B(_15953_), .C(_15954_), .Y(_15961_) );
NAND2X1 NAND2X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_15961_), .B(_15960_), .Y(_15962_) );
NAND3X1 NAND3X1_3678 ( .gnd(gnd), .vdd(vdd), .A(_15959_), .B(_14296_), .C(_15962_), .Y(_15963_) );
NAND3X1 NAND3X1_3679 ( .gnd(gnd), .vdd(vdd), .A(_15736_), .B(_15963_), .C(_15958_), .Y(_15964_) );
NAND3X1 NAND3X1_3680 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_190_), .B(_14296_), .C(_15962_), .Y(_15965_) );
NAND2X1 NAND2X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_15959_), .B(_15956_), .Y(_15966_) );
NAND3X1 NAND3X1_3681 ( .gnd(gnd), .vdd(vdd), .A(_15632_), .B(_15965_), .C(_15966_), .Y(_15967_) );
AOI21X1 AOI21X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_15964_), .B(_15967_), .C(_15735_), .Y(_15969_) );
NAND3X1 NAND3X1_3682 ( .gnd(gnd), .vdd(vdd), .A(_15632_), .B(_15963_), .C(_15958_), .Y(_15970_) );
NAND3X1 NAND3X1_3683 ( .gnd(gnd), .vdd(vdd), .A(_15736_), .B(_15965_), .C(_15966_), .Y(_15971_) );
AOI21X1 AOI21X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_15970_), .B(_15971_), .C(_15734_), .Y(_15972_) );
OAI21X1 OAI21X1_2536 ( .gnd(gnd), .vdd(vdd), .A(_15969_), .B(_15972_), .C(_13867_), .Y(_15973_) );
NAND3X1 NAND3X1_3684 ( .gnd(gnd), .vdd(vdd), .A(_15734_), .B(_15970_), .C(_15971_), .Y(_15974_) );
NAND3X1 NAND3X1_3685 ( .gnd(gnd), .vdd(vdd), .A(_15964_), .B(_15967_), .C(_15735_), .Y(_15975_) );
NAND3X1 NAND3X1_3686 ( .gnd(gnd), .vdd(vdd), .A(_13868_), .B(_15974_), .C(_15975_), .Y(_15976_) );
NAND3X1 NAND3X1_3687 ( .gnd(gnd), .vdd(vdd), .A(_14332_), .B(_15976_), .C(_15973_), .Y(_15977_) );
NAND2X1 NAND2X1_2048 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_206_), .B(_15977_), .Y(_15978_) );
INVX1 INVX1_2202 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_206_), .Y(_15980_) );
NAND3X1 NAND3X1_3688 ( .gnd(gnd), .vdd(vdd), .A(_13867_), .B(_15974_), .C(_15975_), .Y(_15981_) );
OAI21X1 OAI21X1_2537 ( .gnd(gnd), .vdd(vdd), .A(_15969_), .B(_15972_), .C(_13868_), .Y(_15982_) );
NAND2X1 NAND2X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_15981_), .B(_15982_), .Y(_15983_) );
NAND3X1 NAND3X1_3689 ( .gnd(gnd), .vdd(vdd), .A(_15980_), .B(_14332_), .C(_15983_), .Y(_15984_) );
NAND3X1 NAND3X1_3690 ( .gnd(gnd), .vdd(vdd), .A(_15647_), .B(_15984_), .C(_15978_), .Y(_15985_) );
INVX1 INVX1_2203 ( .gnd(gnd), .vdd(vdd), .A(_15647_), .Y(_15986_) );
NAND3X1 NAND3X1_3691 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_206_), .B(_14332_), .C(_15983_), .Y(_15987_) );
NAND2X1 NAND2X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_15980_), .B(_15977_), .Y(_15988_) );
NAND3X1 NAND3X1_3692 ( .gnd(gnd), .vdd(vdd), .A(_15986_), .B(_15987_), .C(_15988_), .Y(_15989_) );
NAND3X1 NAND3X1_3693 ( .gnd(gnd), .vdd(vdd), .A(_15733_), .B(_15985_), .C(_15989_), .Y(_15991_) );
AOI21X1 AOI21X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_15662_), .B(_15659_), .C(_15653_), .Y(_15992_) );
AOI21X1 AOI21X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_15987_), .B(_15988_), .C(_15986_), .Y(_15993_) );
AOI21X1 AOI21X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_15984_), .B(_15978_), .C(_15647_), .Y(_15994_) );
OAI21X1 OAI21X1_2538 ( .gnd(gnd), .vdd(vdd), .A(_15993_), .B(_15994_), .C(_15992_), .Y(_15995_) );
NAND3X1 NAND3X1_3694 ( .gnd(gnd), .vdd(vdd), .A(_13864_), .B(_15991_), .C(_15995_), .Y(_15996_) );
NOR3X1 NOR3X1_469 ( .gnd(gnd), .vdd(vdd), .A(_15993_), .B(_15992_), .C(_15994_), .Y(_15997_) );
AOI21X1 AOI21X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_15985_), .B(_15989_), .C(_15733_), .Y(_15998_) );
OAI21X1 OAI21X1_2539 ( .gnd(gnd), .vdd(vdd), .A(_15997_), .B(_15998_), .C(_16517_), .Y(_15999_) );
NAND3X1 NAND3X1_3695 ( .gnd(gnd), .vdd(vdd), .A(_14369_), .B(_15996_), .C(_15999_), .Y(_16000_) );
NAND2X1 NAND2X1_2051 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_222_), .B(_16000_), .Y(_16002_) );
INVX1 INVX1_2204 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_222_), .Y(_16003_) );
NAND2X1 NAND2X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_15991_), .B(_15995_), .Y(_16004_) );
AOI21X1 AOI21X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_16517_), .B(_16004_), .C(_14370_), .Y(_16005_) );
NAND3X1 NAND3X1_3696 ( .gnd(gnd), .vdd(vdd), .A(_16003_), .B(_15996_), .C(_16005_), .Y(_16006_) );
NAND3X1 NAND3X1_3697 ( .gnd(gnd), .vdd(vdd), .A(_15676_), .B(_16006_), .C(_16002_), .Y(_16007_) );
INVX1 INVX1_2205 ( .gnd(gnd), .vdd(vdd), .A(_15676_), .Y(_16008_) );
NAND3X1 NAND3X1_3698 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_222_), .B(_15996_), .C(_16005_), .Y(_16009_) );
NAND2X1 NAND2X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_16003_), .B(_16000_), .Y(_16010_) );
NAND3X1 NAND3X1_3699 ( .gnd(gnd), .vdd(vdd), .A(_16008_), .B(_16009_), .C(_16010_), .Y(_16011_) );
NAND3X1 NAND3X1_3700 ( .gnd(gnd), .vdd(vdd), .A(_15732_), .B(_16007_), .C(_16011_), .Y(_16013_) );
AOI21X1 AOI21X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_15678_), .B(_15367_), .C(_15681_), .Y(_16014_) );
NAND3X1 NAND3X1_3701 ( .gnd(gnd), .vdd(vdd), .A(_16008_), .B(_16006_), .C(_16002_), .Y(_16015_) );
NAND3X1 NAND3X1_3702 ( .gnd(gnd), .vdd(vdd), .A(_15676_), .B(_16009_), .C(_16010_), .Y(_16016_) );
NAND3X1 NAND3X1_3703 ( .gnd(gnd), .vdd(vdd), .A(_16014_), .B(_16015_), .C(_16016_), .Y(_16017_) );
NAND3X1 NAND3X1_3704 ( .gnd(gnd), .vdd(vdd), .A(_13861_), .B(_16013_), .C(_16017_), .Y(_16018_) );
AOI21X1 AOI21X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_16015_), .B(_16016_), .C(_16014_), .Y(_16019_) );
AOI21X1 AOI21X1_2252 ( .gnd(gnd), .vdd(vdd), .A(_16007_), .B(_16011_), .C(_15732_), .Y(_16020_) );
OAI21X1 OAI21X1_2540 ( .gnd(gnd), .vdd(vdd), .A(_16019_), .B(_16020_), .C(_13860_), .Y(_16021_) );
NAND3X1 NAND3X1_3705 ( .gnd(gnd), .vdd(vdd), .A(_14406_), .B(_16018_), .C(_16021_), .Y(_16022_) );
NAND2X1 NAND2X1_2054 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_238_), .B(_16022_), .Y(_16024_) );
INVX1 INVX1_2206 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_238_), .Y(_16025_) );
NAND2X1 NAND2X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_16013_), .B(_16017_), .Y(_16026_) );
AOI21X1 AOI21X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_13860_), .B(_16026_), .C(_14407_), .Y(_16027_) );
NAND3X1 NAND3X1_3706 ( .gnd(gnd), .vdd(vdd), .A(_16025_), .B(_16018_), .C(_16027_), .Y(_16028_) );
NAND3X1 NAND3X1_3707 ( .gnd(gnd), .vdd(vdd), .A(_15691_), .B(_16028_), .C(_16024_), .Y(_16029_) );
INVX2 INVX2_536 ( .gnd(gnd), .vdd(vdd), .A(_15691_), .Y(_16030_) );
NAND3X1 NAND3X1_3708 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_238_), .B(_16018_), .C(_16027_), .Y(_16031_) );
NAND2X1 NAND2X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_16025_), .B(_16022_), .Y(_16032_) );
NAND3X1 NAND3X1_3709 ( .gnd(gnd), .vdd(vdd), .A(_16030_), .B(_16031_), .C(_16032_), .Y(_16033_) );
NAND3X1 NAND3X1_3710 ( .gnd(gnd), .vdd(vdd), .A(_16029_), .B(_16033_), .C(_15731_), .Y(_16035_) );
AOI21X1 AOI21X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_15706_), .B(_15703_), .C(_15697_), .Y(_16036_) );
AOI21X1 AOI21X1_2255 ( .gnd(gnd), .vdd(vdd), .A(_16031_), .B(_16032_), .C(_16030_), .Y(_16037_) );
AOI21X1 AOI21X1_2256 ( .gnd(gnd), .vdd(vdd), .A(_16028_), .B(_16024_), .C(_15691_), .Y(_16038_) );
OAI21X1 OAI21X1_2541 ( .gnd(gnd), .vdd(vdd), .A(_16037_), .B(_16038_), .C(_16036_), .Y(_16039_) );
NAND3X1 NAND3X1_3711 ( .gnd(gnd), .vdd(vdd), .A(_16767_), .B(_16035_), .C(_16039_), .Y(_16040_) );
NAND3X1 NAND3X1_3712 ( .gnd(gnd), .vdd(vdd), .A(_16030_), .B(_16028_), .C(_16024_), .Y(_16041_) );
NAND3X1 NAND3X1_3713 ( .gnd(gnd), .vdd(vdd), .A(_15691_), .B(_16031_), .C(_16032_), .Y(_16042_) );
AOI21X1 AOI21X1_2257 ( .gnd(gnd), .vdd(vdd), .A(_16041_), .B(_16042_), .C(_16036_), .Y(_16043_) );
AOI21X1 AOI21X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_16029_), .B(_16033_), .C(_15731_), .Y(_16044_) );
OAI21X1 OAI21X1_2542 ( .gnd(gnd), .vdd(vdd), .A(_16043_), .B(_16044_), .C(_16539_), .Y(_16046_) );
NAND3X1 NAND3X1_3714 ( .gnd(gnd), .vdd(vdd), .A(_14441_), .B(_16040_), .C(_16046_), .Y(_16047_) );
NAND2X1 NAND2X1_2057 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_254_), .B(_16047_), .Y(_16048_) );
INVX1 INVX1_2207 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_254_), .Y(_16049_) );
NAND2X1 NAND2X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_16035_), .B(_16039_), .Y(_16050_) );
AOI21X1 AOI21X1_2259 ( .gnd(gnd), .vdd(vdd), .A(_16539_), .B(_16050_), .C(_14442_), .Y(_16051_) );
NAND3X1 NAND3X1_3715 ( .gnd(gnd), .vdd(vdd), .A(_16049_), .B(_16040_), .C(_16051_), .Y(_16052_) );
NAND3X1 NAND3X1_3716 ( .gnd(gnd), .vdd(vdd), .A(_15730_), .B(_16052_), .C(_16048_), .Y(_16053_) );
INVX1 INVX1_2208 ( .gnd(gnd), .vdd(vdd), .A(_16053_), .Y(_16054_) );
AOI21X1 AOI21X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_16052_), .B(_16048_), .C(_15730_), .Y(_16055_) );
OAI21X1 OAI21X1_2543 ( .gnd(gnd), .vdd(vdd), .A(_16054_), .B(_16055_), .C(_15729_), .Y(_16057_) );
INVX1 INVX1_2209 ( .gnd(gnd), .vdd(vdd), .A(_16055_), .Y(_16058_) );
NAND3X1 NAND3X1_3717 ( .gnd(gnd), .vdd(vdd), .A(_15728_), .B(_16053_), .C(_16058_), .Y(_16059_) );
NAND2X1 NAND2X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_16057_), .B(_16059_), .Y(module_3_H_22_) );
OAI21X1 OAI21X1_2544 ( .gnd(gnd), .vdd(vdd), .A(_15728_), .B(_16055_), .C(_16053_), .Y(_16060_) );
AOI21X1 AOI21X1_2261 ( .gnd(gnd), .vdd(vdd), .A(_16040_), .B(_16051_), .C(_16049_), .Y(_16061_) );
INVX1 INVX1_2210 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_255_), .Y(_16062_) );
OAI21X1 OAI21X1_2545 ( .gnd(gnd), .vdd(vdd), .A(_16036_), .B(_16038_), .C(_16029_), .Y(_16063_) );
INVX1 INVX1_2211 ( .gnd(gnd), .vdd(vdd), .A(_16063_), .Y(_16064_) );
NAND2X1 NAND2X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_16007_), .B(_16013_), .Y(_16065_) );
OAI21X1 OAI21X1_2546 ( .gnd(gnd), .vdd(vdd), .A(_15994_), .B(_15992_), .C(_15985_), .Y(_16067_) );
NAND2X1 NAND2X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_15970_), .B(_15974_), .Y(_16068_) );
NAND2X1 NAND2X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_15949_), .B(_15953_), .Y(_16069_) );
INVX1 INVX1_2212 ( .gnd(gnd), .vdd(vdd), .A(_16069_), .Y(_16070_) );
NAND2X1 NAND2X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_15928_), .B(_15932_), .Y(_16071_) );
NAND2X1 NAND2X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .B(_15906_), .Y(_16072_) );
NAND2X1 NAND2X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_15884_), .B(_15889_), .Y(_16073_) );
INVX1 INVX1_2213 ( .gnd(gnd), .vdd(vdd), .A(_16073_), .Y(_16074_) );
INVX1 INVX1_2214 ( .gnd(gnd), .vdd(vdd), .A(_15879_), .Y(_16075_) );
NOR2X1 NOR2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_16673_), .B(_16675_), .Y(_16076_) );
NAND2X1 NAND2X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_15856_), .B(_15861_), .Y(_16078_) );
INVX1 INVX1_2215 ( .gnd(gnd), .vdd(vdd), .A(_16078_), .Y(_16079_) );
OAI21X1 OAI21X1_2547 ( .gnd(gnd), .vdd(vdd), .A(_15842_), .B(_15840_), .C(_15834_), .Y(_16080_) );
INVX1 INVX1_2216 ( .gnd(gnd), .vdd(vdd), .A(_16655_), .Y(_16081_) );
NAND2X1 NAND2X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_15812_), .B(_15817_), .Y(_16082_) );
INVX1 INVX1_2217 ( .gnd(gnd), .vdd(vdd), .A(_16082_), .Y(_16083_) );
NAND2X1 NAND2X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_15790_), .B(_15795_), .Y(_16084_) );
INVX1 INVX1_2218 ( .gnd(gnd), .vdd(vdd), .A(_14693_), .Y(_16085_) );
XNOR2X1 XNOR2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_15785_), .B(_16085_), .Y(_16086_) );
INVX1 INVX1_2219 ( .gnd(gnd), .vdd(vdd), .A(_16086_), .Y(_16087_) );
INVX1 INVX1_2220 ( .gnd(gnd), .vdd(vdd), .A(_15752_), .Y(_16089_) );
NAND2X1 NAND2X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_15772_), .B(_15775_), .Y(_16090_) );
OAI21X1 OAI21X1_2548 ( .gnd(gnd), .vdd(vdd), .A(_16090_), .B(_16089_), .C(_15772_), .Y(_16091_) );
INVX1 INVX1_2221 ( .gnd(gnd), .vdd(vdd), .A(_16091_), .Y(_16092_) );
INVX1 INVX1_2222 ( .gnd(gnd), .vdd(vdd), .A(_15767_), .Y(_16093_) );
OAI21X1 OAI21X1_2549 ( .gnd(gnd), .vdd(vdd), .A(_15423_), .B(_15428_), .C(_15763_), .Y(_16094_) );
OAI21X1 OAI21X1_2550 ( .gnd(gnd), .vdd(vdd), .A(_15417_), .B(_15762_), .C(_16094_), .Y(_16095_) );
INVX1 INVX1_2223 ( .gnd(gnd), .vdd(vdd), .A(_16095_), .Y(_16096_) );
OAI21X1 OAI21X1_2551 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_12_), .B(module_3_W_13_), .C(module_3_W_14_), .Y(_16097_) );
XOR2X1 XOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_11_), .B(module_3_W_15_), .Y(_16098_) );
XNOR2X1 XNOR2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_16098_), .B(_16097_), .Y(_16100_) );
XOR2X1 XOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_16590_), .B(module_3_W_31_), .Y(_16101_) );
XNOR2X1 XNOR2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_16101_), .B(_16100_), .Y(_16102_) );
XOR2X1 XOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_15760_), .B(_16102_), .Y(_16103_) );
XNOR2X1 XNOR2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_16103_), .B(_14489_), .Y(_16104_) );
XNOR2X1 XNOR2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_14657_), .B(bloque_datos[15]), .Y(_16105_) );
XNOR2X1 XNOR2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_16104_), .B(_16105_), .Y(_16106_) );
NOR2X1 NOR2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_16096_), .B(_16106_), .Y(_16107_) );
NAND2X1 NAND2X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_16096_), .B(_16106_), .Y(_16108_) );
INVX1 INVX1_2224 ( .gnd(gnd), .vdd(vdd), .A(_16108_), .Y(_16109_) );
OR2X2 OR2X2_365 ( .gnd(gnd), .vdd(vdd), .A(_16109_), .B(_16107_), .Y(_16111_) );
NOR2X1 NOR2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_16093_), .B(_16111_), .Y(_16112_) );
INVX1 INVX1_2225 ( .gnd(gnd), .vdd(vdd), .A(_16112_), .Y(_16113_) );
OAI21X1 OAI21X1_2552 ( .gnd(gnd), .vdd(vdd), .A(_16109_), .B(_16107_), .C(_16093_), .Y(_16114_) );
XNOR2X1 XNOR2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_14671_), .B(_14495_), .Y(_16115_) );
INVX1 INVX1_2226 ( .gnd(gnd), .vdd(vdd), .A(_16115_), .Y(_16116_) );
NAND3X1 NAND3X1_3718 ( .gnd(gnd), .vdd(vdd), .A(_16114_), .B(_16116_), .C(_16113_), .Y(_16117_) );
AOI21X1 AOI21X1_2262 ( .gnd(gnd), .vdd(vdd), .A(_16114_), .B(_16113_), .C(_16116_), .Y(_16118_) );
INVX1 INVX1_2227 ( .gnd(gnd), .vdd(vdd), .A(_16118_), .Y(_16119_) );
NAND2X1 NAND2X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_16117_), .B(_16119_), .Y(_16120_) );
NOR2X1 NOR2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf3_), .B(_16120_), .Y(_16122_) );
AND2X2 AND2X2_348 ( .gnd(gnd), .vdd(vdd), .A(_16120_), .B(bloque_datos_31_bF_buf2_), .Y(_16123_) );
NOR2X1 NOR2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_16122_), .B(_16123_), .Y(_16124_) );
NAND2X1 NAND2X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_16092_), .B(_16124_), .Y(_16125_) );
OAI21X1 OAI21X1_2553 ( .gnd(gnd), .vdd(vdd), .A(_16123_), .B(_16122_), .C(_16091_), .Y(_16126_) );
XOR2X1 XOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_14510_), .B(bloque_datos_47_bF_buf3_), .Y(_16127_) );
NAND3X1 NAND3X1_3719 ( .gnd(gnd), .vdd(vdd), .A(_16126_), .B(_16127_), .C(_16125_), .Y(_16128_) );
AND2X2 AND2X2_349 ( .gnd(gnd), .vdd(vdd), .A(_16124_), .B(_16092_), .Y(_16129_) );
NOR2X1 NOR2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_16092_), .B(_16124_), .Y(_16130_) );
INVX1 INVX1_2228 ( .gnd(gnd), .vdd(vdd), .A(_16127_), .Y(_16131_) );
OAI21X1 OAI21X1_2554 ( .gnd(gnd), .vdd(vdd), .A(_16129_), .B(_16130_), .C(_16131_), .Y(_16133_) );
AOI21X1 AOI21X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_16128_), .B(_16133_), .C(_16087_), .Y(_16134_) );
INVX1 INVX1_2229 ( .gnd(gnd), .vdd(vdd), .A(_16134_), .Y(_16135_) );
NAND3X1 NAND3X1_3720 ( .gnd(gnd), .vdd(vdd), .A(_16087_), .B(_16128_), .C(_16133_), .Y(_16136_) );
NAND3X1 NAND3X1_3721 ( .gnd(gnd), .vdd(vdd), .A(_16084_), .B(_16136_), .C(_16135_), .Y(_16137_) );
INVX1 INVX1_2230 ( .gnd(gnd), .vdd(vdd), .A(_16084_), .Y(_16138_) );
INVX1 INVX1_2231 ( .gnd(gnd), .vdd(vdd), .A(_16136_), .Y(_16139_) );
OAI21X1 OAI21X1_2555 ( .gnd(gnd), .vdd(vdd), .A(_16139_), .B(_16134_), .C(_16138_), .Y(_16140_) );
OAI21X1 OAI21X1_2556 ( .gnd(gnd), .vdd(vdd), .A(_14521_), .B(_14518_), .C(_16811_), .Y(_16141_) );
NAND2X1 NAND2X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_16640_), .B(_14645_), .Y(_16142_) );
NAND2X1 NAND2X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_16141_), .B(_16142_), .Y(_16144_) );
AOI21X1 AOI21X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_16140_), .B(_16137_), .C(_16144_), .Y(_16145_) );
NAND3X1 NAND3X1_3722 ( .gnd(gnd), .vdd(vdd), .A(_16138_), .B(_16136_), .C(_16135_), .Y(_16146_) );
OAI21X1 OAI21X1_2557 ( .gnd(gnd), .vdd(vdd), .A(_16139_), .B(_16134_), .C(_16084_), .Y(_16147_) );
AOI22X1 AOI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_16141_), .B(_16142_), .C(_16146_), .D(_16147_), .Y(_16148_) );
NOR2X1 NOR2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_16145_), .B(_16148_), .Y(_16149_) );
XNOR2X1 XNOR2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_15807_), .B(bloque_datos[63]), .Y(_16150_) );
AND2X2 AND2X2_350 ( .gnd(gnd), .vdd(vdd), .A(_16149_), .B(_16150_), .Y(_16151_) );
NOR2X1 NOR2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_16150_), .B(_16149_), .Y(_16152_) );
OAI21X1 OAI21X1_2558 ( .gnd(gnd), .vdd(vdd), .A(_16151_), .B(_16152_), .C(_16083_), .Y(_16153_) );
NAND2X1 NAND2X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_16150_), .B(_16149_), .Y(_16155_) );
OR2X2 OR2X2_366 ( .gnd(gnd), .vdd(vdd), .A(_16149_), .B(_16150_), .Y(_16156_) );
NAND3X1 NAND3X1_3723 ( .gnd(gnd), .vdd(vdd), .A(_16082_), .B(_16155_), .C(_16156_), .Y(_16157_) );
NAND3X1 NAND3X1_3724 ( .gnd(gnd), .vdd(vdd), .A(_16081_), .B(_16153_), .C(_16157_), .Y(_16158_) );
NAND3X1 NAND3X1_3725 ( .gnd(gnd), .vdd(vdd), .A(_16083_), .B(_16155_), .C(_16156_), .Y(_16159_) );
OAI21X1 OAI21X1_2559 ( .gnd(gnd), .vdd(vdd), .A(_16151_), .B(_16152_), .C(_16082_), .Y(_16160_) );
NAND3X1 NAND3X1_3726 ( .gnd(gnd), .vdd(vdd), .A(_16655_), .B(_16160_), .C(_16159_), .Y(_16161_) );
NAND2X1 NAND2X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_16158_), .B(_16161_), .Y(_16162_) );
XOR2X1 XOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_14643_), .B(bloque_datos_79_bF_buf3_), .Y(_16163_) );
NOR2X1 NOR2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_15829_), .B(_16163_), .Y(_16164_) );
INVX1 INVX1_2232 ( .gnd(gnd), .vdd(vdd), .A(_16164_), .Y(_16166_) );
NAND2X1 NAND2X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_15829_), .B(_16163_), .Y(_16167_) );
NAND2X1 NAND2X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_16167_), .B(_16166_), .Y(_16168_) );
NAND2X1 NAND2X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_16168_), .B(_16162_), .Y(_16169_) );
OR2X2 OR2X2_367 ( .gnd(gnd), .vdd(vdd), .A(_16162_), .B(_16168_), .Y(_16170_) );
NAND3X1 NAND3X1_3727 ( .gnd(gnd), .vdd(vdd), .A(_16080_), .B(_16169_), .C(_16170_), .Y(_16171_) );
INVX1 INVX1_2233 ( .gnd(gnd), .vdd(vdd), .A(_16080_), .Y(_16172_) );
AND2X2 AND2X2_351 ( .gnd(gnd), .vdd(vdd), .A(_16162_), .B(_16168_), .Y(_16173_) );
NOR2X1 NOR2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_16168_), .B(_16162_), .Y(_16174_) );
OAI21X1 OAI21X1_2560 ( .gnd(gnd), .vdd(vdd), .A(_16173_), .B(_16174_), .C(_16172_), .Y(_16175_) );
NOR2X1 NOR2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_16661_), .B(_16663_), .Y(_16177_) );
XNOR2X1 XNOR2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_14641_), .B(_16177_), .Y(_16178_) );
INVX1 INVX1_2234 ( .gnd(gnd), .vdd(vdd), .A(_16178_), .Y(_16179_) );
AOI21X1 AOI21X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_16175_), .B(_16171_), .C(_16179_), .Y(_16180_) );
NAND3X1 NAND3X1_3728 ( .gnd(gnd), .vdd(vdd), .A(_16172_), .B(_16169_), .C(_16170_), .Y(_16181_) );
OAI21X1 OAI21X1_2561 ( .gnd(gnd), .vdd(vdd), .A(_16173_), .B(_16174_), .C(_16080_), .Y(_16182_) );
AOI21X1 AOI21X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_16182_), .B(_16181_), .C(_16178_), .Y(_16183_) );
NOR2X1 NOR2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_16180_), .B(_16183_), .Y(_16184_) );
NAND2X1 NAND2X1_2080 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf3_), .B(_15851_), .Y(_16185_) );
NOR2X1 NOR2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf2_), .B(_15851_), .Y(_16186_) );
INVX1 INVX1_2235 ( .gnd(gnd), .vdd(vdd), .A(_16186_), .Y(_16188_) );
NAND2X1 NAND2X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_16185_), .B(_16188_), .Y(_16189_) );
NAND2X1 NAND2X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_16189_), .B(_16184_), .Y(_16190_) );
OR2X2 OR2X2_368 ( .gnd(gnd), .vdd(vdd), .A(_16184_), .B(_16189_), .Y(_16191_) );
NAND3X1 NAND3X1_3729 ( .gnd(gnd), .vdd(vdd), .A(_16079_), .B(_16190_), .C(_16191_), .Y(_16192_) );
AND2X2 AND2X2_352 ( .gnd(gnd), .vdd(vdd), .A(_16184_), .B(_16189_), .Y(_16193_) );
NOR2X1 NOR2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_16189_), .B(_16184_), .Y(_16194_) );
OAI21X1 OAI21X1_2562 ( .gnd(gnd), .vdd(vdd), .A(_16193_), .B(_16194_), .C(_16078_), .Y(_16195_) );
AOI21X1 AOI21X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_16195_), .B(_16192_), .C(_16076_), .Y(_16196_) );
INVX1 INVX1_2236 ( .gnd(gnd), .vdd(vdd), .A(_16076_), .Y(_16197_) );
OAI21X1 OAI21X1_2563 ( .gnd(gnd), .vdd(vdd), .A(_16193_), .B(_16194_), .C(_16079_), .Y(_16199_) );
NAND3X1 NAND3X1_3730 ( .gnd(gnd), .vdd(vdd), .A(_16078_), .B(_16190_), .C(_16191_), .Y(_16200_) );
AOI21X1 AOI21X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_16199_), .B(_16200_), .C(_16197_), .Y(_16201_) );
OAI21X1 OAI21X1_2564 ( .gnd(gnd), .vdd(vdd), .A(_16196_), .B(_16201_), .C(_16075_), .Y(_16202_) );
NAND3X1 NAND3X1_3731 ( .gnd(gnd), .vdd(vdd), .A(_16197_), .B(_16199_), .C(_16200_), .Y(_16203_) );
NAND3X1 NAND3X1_3732 ( .gnd(gnd), .vdd(vdd), .A(_16076_), .B(_16195_), .C(_16192_), .Y(_16204_) );
NAND3X1 NAND3X1_3733 ( .gnd(gnd), .vdd(vdd), .A(_15879_), .B(_16203_), .C(_16204_), .Y(_16205_) );
NAND2X1 NAND2X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_16205_), .B(_16202_), .Y(_16206_) );
AOI21X1 AOI21X1_2269 ( .gnd(gnd), .vdd(vdd), .A(_16074_), .B(_16206_), .C(_14554_), .Y(_16207_) );
OAI21X1 OAI21X1_2565 ( .gnd(gnd), .vdd(vdd), .A(_16074_), .B(_16206_), .C(_16207_), .Y(_16208_) );
XOR2X1 XOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_14810_), .B(module_3_W_143_), .Y(_16210_) );
XOR2X1 XOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_16208_), .B(_16210_), .Y(_16211_) );
XOR2X1 XOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_16211_), .B(_15894_), .Y(_16212_) );
NAND2X1 NAND2X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_16072_), .B(_16212_), .Y(_16213_) );
INVX1 INVX1_2237 ( .gnd(gnd), .vdd(vdd), .A(_16072_), .Y(_16214_) );
XNOR2X1 XNOR2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_16211_), .B(_15894_), .Y(_16215_) );
AOI21X1 AOI21X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_16214_), .B(_16215_), .C(_14808_), .Y(_16216_) );
XNOR2X1 XNOR2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_16698_), .B(module_3_W_159_), .Y(_16217_) );
NAND3X1 NAND3X1_3734 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_16217_), .C(_16216_), .Y(_16218_) );
NOR2X1 NOR2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_16214_), .B(_16215_), .Y(_16219_) );
OAI21X1 OAI21X1_2566 ( .gnd(gnd), .vdd(vdd), .A(_16212_), .B(_16072_), .C(_14563_), .Y(_16221_) );
INVX1 INVX1_2238 ( .gnd(gnd), .vdd(vdd), .A(_16217_), .Y(_16222_) );
OAI21X1 OAI21X1_2567 ( .gnd(gnd), .vdd(vdd), .A(_16221_), .B(_16219_), .C(_16222_), .Y(_16223_) );
NAND2X1 NAND2X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_16218_), .B(_16223_), .Y(_16224_) );
XOR2X1 XOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_16224_), .B(_15917_), .Y(_16225_) );
NAND2X1 NAND2X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_16071_), .B(_16225_), .Y(_16226_) );
INVX1 INVX1_2239 ( .gnd(gnd), .vdd(vdd), .A(_16071_), .Y(_16227_) );
XNOR2X1 XNOR2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_16224_), .B(_15917_), .Y(_16228_) );
AOI21X1 AOI21X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_16227_), .B(_16228_), .C(_14576_), .Y(_16229_) );
XOR2X1 XOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_16709_), .B(module_3_W_175_), .Y(_16230_) );
NAND3X1 NAND3X1_3735 ( .gnd(gnd), .vdd(vdd), .A(_16226_), .B(_16230_), .C(_16229_), .Y(_16232_) );
NOR2X1 NOR2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_16227_), .B(_16228_), .Y(_16233_) );
OAI21X1 OAI21X1_2568 ( .gnd(gnd), .vdd(vdd), .A(_16225_), .B(_16071_), .C(_14637_), .Y(_16234_) );
INVX1 INVX1_2240 ( .gnd(gnd), .vdd(vdd), .A(_16230_), .Y(_16235_) );
OAI21X1 OAI21X1_2569 ( .gnd(gnd), .vdd(vdd), .A(_16234_), .B(_16233_), .C(_16235_), .Y(_16236_) );
NAND2X1 NAND2X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_16232_), .B(_16236_), .Y(_16237_) );
XNOR2X1 XNOR2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_16237_), .B(_15937_), .Y(_16238_) );
NAND2X1 NAND2X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_16070_), .B(_16238_), .Y(_16239_) );
XOR2X1 XOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_16237_), .B(_15937_), .Y(_16240_) );
AOI21X1 AOI21X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_16069_), .B(_16240_), .C(_14586_), .Y(_16241_) );
AND2X2 AND2X2_353 ( .gnd(gnd), .vdd(vdd), .A(_13291_), .B(module_3_W_191_), .Y(_16243_) );
NOR2X1 NOR2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_191_), .B(_13291_), .Y(_16244_) );
NOR2X1 NOR2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_16244_), .B(_16243_), .Y(_16245_) );
NAND3X1 NAND3X1_3736 ( .gnd(gnd), .vdd(vdd), .A(_16239_), .B(_16245_), .C(_16241_), .Y(_16246_) );
NOR2X1 NOR2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_16069_), .B(_16240_), .Y(_16247_) );
OAI21X1 OAI21X1_2570 ( .gnd(gnd), .vdd(vdd), .A(_16238_), .B(_16070_), .C(_14633_), .Y(_16248_) );
OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_16243_), .B(_16244_), .C(_16248_), .D(_16247_), .Y(_16249_) );
NAND2X1 NAND2X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_16246_), .B(_16249_), .Y(_16250_) );
XOR2X1 XOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_16250_), .B(_15958_), .Y(_16251_) );
NAND2X1 NAND2X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_16068_), .B(_16251_), .Y(_16252_) );
INVX1 INVX1_2241 ( .gnd(gnd), .vdd(vdd), .A(_16068_), .Y(_16254_) );
XNOR2X1 XNOR2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_16250_), .B(_15958_), .Y(_16255_) );
AOI21X1 AOI21X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_16254_), .B(_16255_), .C(_14872_), .Y(_16256_) );
OAI21X1 OAI21X1_2571 ( .gnd(gnd), .vdd(vdd), .A(_16730_), .B(_16733_), .C(module_3_W_207_), .Y(_16257_) );
INVX1 INVX1_2242 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_207_), .Y(_16258_) );
NAND3X1 NAND3X1_3737 ( .gnd(gnd), .vdd(vdd), .A(_16258_), .B(_16732_), .C(_16737_), .Y(_16259_) );
NAND2X1 NAND2X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_16259_), .B(_16257_), .Y(_16260_) );
INVX1 INVX1_2243 ( .gnd(gnd), .vdd(vdd), .A(_16260_), .Y(_16261_) );
NAND3X1 NAND3X1_3738 ( .gnd(gnd), .vdd(vdd), .A(_16252_), .B(_16261_), .C(_16256_), .Y(_16262_) );
NOR2X1 NOR2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_16254_), .B(_16255_), .Y(_16263_) );
OAI21X1 OAI21X1_2572 ( .gnd(gnd), .vdd(vdd), .A(_16251_), .B(_16068_), .C(_14595_), .Y(_16265_) );
OAI21X1 OAI21X1_2573 ( .gnd(gnd), .vdd(vdd), .A(_16265_), .B(_16263_), .C(_16260_), .Y(_16266_) );
NAND2X1 NAND2X1_2092 ( .gnd(gnd), .vdd(vdd), .A(_16262_), .B(_16266_), .Y(_16267_) );
XOR2X1 XOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_16267_), .B(_15978_), .Y(_16268_) );
XNOR2X1 XNOR2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_16268_), .B(_16067_), .Y(_16269_) );
OAI21X1 OAI21X1_2574 ( .gnd(gnd), .vdd(vdd), .A(_16745_), .B(_16748_), .C(module_3_W_223_), .Y(_16270_) );
INVX1 INVX1_2244 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_223_), .Y(_16271_) );
NAND2X1 NAND2X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_16271_), .B(_16750_), .Y(_16272_) );
NAND2X1 NAND2X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_16270_), .B(_16272_), .Y(_16273_) );
NOR3X1 NOR3X1_470 ( .gnd(gnd), .vdd(vdd), .A(_16273_), .B(_14606_), .C(_16269_), .Y(_16274_) );
XOR2X1 XOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_16268_), .B(_16067_), .Y(_16276_) );
AND2X2 AND2X2_354 ( .gnd(gnd), .vdd(vdd), .A(_16272_), .B(_16270_), .Y(_16277_) );
AOI21X1 AOI21X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_14885_), .B(_16276_), .C(_16277_), .Y(_16278_) );
OAI21X1 OAI21X1_2575 ( .gnd(gnd), .vdd(vdd), .A(_16274_), .B(_16278_), .C(_16002_), .Y(_16279_) );
INVX1 INVX1_2245 ( .gnd(gnd), .vdd(vdd), .A(_16002_), .Y(_16280_) );
NAND3X1 NAND3X1_3739 ( .gnd(gnd), .vdd(vdd), .A(_14885_), .B(_16276_), .C(_16277_), .Y(_16281_) );
OAI21X1 OAI21X1_2576 ( .gnd(gnd), .vdd(vdd), .A(_16269_), .B(_14606_), .C(_16273_), .Y(_16282_) );
NAND3X1 NAND3X1_3740 ( .gnd(gnd), .vdd(vdd), .A(_16280_), .B(_16281_), .C(_16282_), .Y(_16283_) );
AND2X2 AND2X2_355 ( .gnd(gnd), .vdd(vdd), .A(_16279_), .B(_16283_), .Y(_16284_) );
NAND2X1 NAND2X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_16065_), .B(_16284_), .Y(_16285_) );
INVX1 INVX1_2246 ( .gnd(gnd), .vdd(vdd), .A(_16065_), .Y(_16287_) );
NAND2X1 NAND2X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_16283_), .B(_16279_), .Y(_16288_) );
AOI21X1 AOI21X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_16288_), .B(_16287_), .C(_14616_), .Y(_16289_) );
OAI21X1 OAI21X1_2577 ( .gnd(gnd), .vdd(vdd), .A(_16761_), .B(_16756_), .C(module_3_W_239_), .Y(_16290_) );
INVX1 INVX1_2247 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_239_), .Y(_16291_) );
NAND3X1 NAND3X1_3741 ( .gnd(gnd), .vdd(vdd), .A(_16291_), .B(_16755_), .C(_16760_), .Y(_16292_) );
AND2X2 AND2X2_356 ( .gnd(gnd), .vdd(vdd), .A(_16290_), .B(_16292_), .Y(_16293_) );
NAND3X1 NAND3X1_3742 ( .gnd(gnd), .vdd(vdd), .A(_16285_), .B(_16289_), .C(_16293_), .Y(_16294_) );
NOR2X1 NOR2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_16288_), .B(_16287_), .Y(_16295_) );
OAI21X1 OAI21X1_2578 ( .gnd(gnd), .vdd(vdd), .A(_16284_), .B(_16065_), .C(_14629_), .Y(_16296_) );
NAND2X1 NAND2X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_16292_), .B(_16290_), .Y(_16298_) );
OAI21X1 OAI21X1_2579 ( .gnd(gnd), .vdd(vdd), .A(_16296_), .B(_16295_), .C(_16298_), .Y(_16299_) );
NAND2X1 NAND2X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_16299_), .B(_16294_), .Y(_16300_) );
XNOR2X1 XNOR2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_16300_), .B(_16024_), .Y(_16301_) );
NOR2X1 NOR2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_16064_), .B(_16301_), .Y(_16302_) );
XOR2X1 XOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_16300_), .B(_16024_), .Y(_16303_) );
OAI21X1 OAI21X1_2580 ( .gnd(gnd), .vdd(vdd), .A(_16303_), .B(_16063_), .C(_14628_), .Y(_16304_) );
OAI21X1 OAI21X1_2581 ( .gnd(gnd), .vdd(vdd), .A(_16304_), .B(_16302_), .C(_16062_), .Y(_16305_) );
OAI21X1 OAI21X1_2582 ( .gnd(gnd), .vdd(vdd), .A(_16043_), .B(_16037_), .C(_16303_), .Y(_16306_) );
AOI21X1 AOI21X1_2276 ( .gnd(gnd), .vdd(vdd), .A(_16064_), .B(_16301_), .C(_14627_), .Y(_16307_) );
NAND3X1 NAND3X1_3743 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_255_), .B(_16306_), .C(_16307_), .Y(_16309_) );
NAND3X1 NAND3X1_3744 ( .gnd(gnd), .vdd(vdd), .A(_16061_), .B(_16309_), .C(_16305_), .Y(_16310_) );
NAND3X1 NAND3X1_3745 ( .gnd(gnd), .vdd(vdd), .A(_16062_), .B(_16306_), .C(_16307_), .Y(_16311_) );
OAI21X1 OAI21X1_2583 ( .gnd(gnd), .vdd(vdd), .A(_16304_), .B(_16302_), .C(module_3_W_255_), .Y(_16312_) );
NAND3X1 NAND3X1_3746 ( .gnd(gnd), .vdd(vdd), .A(_16048_), .B(_16311_), .C(_16312_), .Y(_16313_) );
NAND2X1 NAND2X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_16313_), .B(_16310_), .Y(_16314_) );
XNOR2X1 XNOR2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_16060_), .B(_16314_), .Y(module_3_H_23_) );
INVX1 INVX1_2248 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_241_), .Y(_14864_) );
AND2X2 AND2X2_357 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_0_), .B(module_3_W_16_), .Y(_14875_) );
NOR2X1 NOR2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_0_), .B(module_3_W_16_), .Y(_14886_) );
OAI21X1 OAI21X1_2584 ( .gnd(gnd), .vdd(vdd), .A(_14875_), .B(_14886_), .C(bloque_datos[0]), .Y(_14897_) );
INVX1 INVX1_2249 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(_14908_) );
NOR2X1 NOR2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_14886_), .B(_14875_), .Y(_14919_) );
NAND2X1 NAND2X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .B(_14919_), .Y(_14930_) );
NAND2X1 NAND2X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .B(_14930_), .Y(_14941_) );
NAND2X1 NAND2X1_2102 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf3_), .B(_14941_), .Y(_14952_) );
OR2X2 OR2X2_369 ( .gnd(gnd), .vdd(vdd), .A(_14941_), .B(bloque_datos_16_bF_buf2_), .Y(_14963_) );
NAND2X1 NAND2X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_14952_), .B(_14963_), .Y(_14972_) );
NAND2X1 NAND2X1_2104 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf1_), .B(_14972_), .Y(_14981_) );
OR2X2 OR2X2_370 ( .gnd(gnd), .vdd(vdd), .A(_14972_), .B(bloque_datos_32_bF_buf0_), .Y(_14991_) );
NAND2X1 NAND2X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_14981_), .B(_14991_), .Y(_15002_) );
NAND2X1 NAND2X1_2106 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_48_bF_buf1_), .B(_15002_), .Y(_15013_) );
OR2X2 OR2X2_371 ( .gnd(gnd), .vdd(vdd), .A(_15002_), .B(bloque_datos_48_bF_buf0_), .Y(_15024_) );
NAND2X1 NAND2X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_15013_), .B(_15024_), .Y(_15035_) );
NAND2X1 NAND2X1_2108 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_64_bF_buf1_), .B(_15035_), .Y(_15046_) );
OR2X2 OR2X2_372 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(bloque_datos_64_bF_buf0_), .Y(_15057_) );
NAND2X1 NAND2X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_15046_), .B(_15057_), .Y(_15068_) );
NAND2X1 NAND2X1_2110 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf5_), .B(_15068_), .Y(_15079_) );
OR2X2 OR2X2_373 ( .gnd(gnd), .vdd(vdd), .A(_15068_), .B(bloque_datos_80_bF_buf4_), .Y(_15090_) );
NAND2X1 NAND2X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_15079_), .B(_15090_), .Y(_15101_) );
NAND2X1 NAND2X1_2112 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_128_), .B(_15101_), .Y(_15112_) );
OR2X2 OR2X2_374 ( .gnd(gnd), .vdd(vdd), .A(_15101_), .B(module_3_W_128_), .Y(_15123_) );
NAND2X1 NAND2X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_15112_), .B(_15123_), .Y(_15134_) );
NAND2X1 NAND2X1_2114 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_144_), .B(_15134_), .Y(_15145_) );
OR2X2 OR2X2_375 ( .gnd(gnd), .vdd(vdd), .A(_15134_), .B(module_3_W_144_), .Y(_15156_) );
NAND2X1 NAND2X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_15145_), .B(_15156_), .Y(_15167_) );
NAND2X1 NAND2X1_2116 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_160_), .B(_15167_), .Y(_15178_) );
OR2X2 OR2X2_376 ( .gnd(gnd), .vdd(vdd), .A(_15167_), .B(module_3_W_160_), .Y(_15189_) );
NAND2X1 NAND2X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_15178_), .B(_15189_), .Y(_15200_) );
NAND2X1 NAND2X1_2118 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_176_), .B(_15200_), .Y(_15211_) );
OR2X2 OR2X2_377 ( .gnd(gnd), .vdd(vdd), .A(_15200_), .B(module_3_W_176_), .Y(_15222_) );
NAND2X1 NAND2X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_15211_), .B(_15222_), .Y(_15233_) );
NAND2X1 NAND2X1_2120 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_192_), .B(_15233_), .Y(_15244_) );
OR2X2 OR2X2_378 ( .gnd(gnd), .vdd(vdd), .A(_15233_), .B(module_3_W_192_), .Y(_15255_) );
NAND2X1 NAND2X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_15244_), .B(_15255_), .Y(_15266_) );
NAND2X1 NAND2X1_2122 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_208_), .B(_15266_), .Y(_15277_) );
OR2X2 OR2X2_379 ( .gnd(gnd), .vdd(vdd), .A(_15266_), .B(module_3_W_208_), .Y(_15288_) );
NAND2X1 NAND2X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_15277_), .B(_15288_), .Y(_15299_) );
INVX2 INVX2_537 ( .gnd(gnd), .vdd(vdd), .A(_15299_), .Y(_15310_) );
NOR2X1 NOR2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_224_), .B(_15310_), .Y(_15321_) );
INVX1 INVX1_2250 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_225_), .Y(_15332_) );
INVX2 INVX2_538 ( .gnd(gnd), .vdd(vdd), .A(_15266_), .Y(_15343_) );
NOR2X1 NOR2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_208_), .B(_15343_), .Y(_15354_) );
INVX2 INVX2_539 ( .gnd(gnd), .vdd(vdd), .A(_15233_), .Y(_15364_) );
NOR2X1 NOR2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_192_), .B(_15364_), .Y(_15375_) );
INVX1 INVX1_2251 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_193_), .Y(_15386_) );
INVX2 INVX2_540 ( .gnd(gnd), .vdd(vdd), .A(_15200_), .Y(_15397_) );
NOR2X1 NOR2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_176_), .B(_15397_), .Y(_15408_) );
INVX2 INVX2_541 ( .gnd(gnd), .vdd(vdd), .A(_15167_), .Y(_15419_) );
NOR2X1 NOR2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_160_), .B(_15419_), .Y(_15430_) );
INVX1 INVX1_2252 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_161_), .Y(_15441_) );
INVX2 INVX2_542 ( .gnd(gnd), .vdd(vdd), .A(_15134_), .Y(_15452_) );
NOR2X1 NOR2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_144_), .B(_15452_), .Y(_15463_) );
INVX1 INVX1_2253 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_145_), .Y(_15474_) );
INVX2 INVX2_543 ( .gnd(gnd), .vdd(vdd), .A(_15101_), .Y(_15485_) );
NOR2X1 NOR2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_128_), .B(_15485_), .Y(_15496_) );
INVX2 INVX2_544 ( .gnd(gnd), .vdd(vdd), .A(_15068_), .Y(_15507_) );
NOR2X1 NOR2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf3_), .B(_15507_), .Y(_15518_) );
AOI21X1 AOI21X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_15013_), .B(_15024_), .C(bloque_datos_64_bF_buf4_), .Y(_15529_) );
AOI21X1 AOI21X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_14981_), .B(_14991_), .C(bloque_datos_48_bF_buf4_), .Y(_15540_) );
INVX1 INVX1_2254 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_49_bF_buf3_), .Y(_15551_) );
AOI21X1 AOI21X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_14952_), .B(_14963_), .C(bloque_datos_32_bF_buf4_), .Y(_15562_) );
INVX1 INVX1_2255 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf0_), .Y(_15573_) );
AOI21X1 AOI21X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .B(_14930_), .C(bloque_datos_16_bF_buf1_), .Y(_15584_) );
OAI21X1 OAI21X1_2585 ( .gnd(gnd), .vdd(vdd), .A(_14875_), .B(_14886_), .C(_14908_), .Y(_15595_) );
INVX1 INVX1_2256 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(_15606_) );
INVX2 INVX2_545 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_0_), .Y(_15617_) );
NOR2X1 NOR2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_16_), .B(_15617_), .Y(_15628_) );
NAND2X1 NAND2X1_2124 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_0_), .B(module_3_W_1_), .Y(_15639_) );
OR2X2 OR2X2_380 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_0_), .B(module_3_W_1_), .Y(_15650_) );
AOI21X1 AOI21X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_15639_), .B(_15650_), .C(module_3_W_17_), .Y(_15661_) );
INVX1 INVX1_2257 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_17_), .Y(_15672_) );
AND2X2 AND2X2_358 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_0_), .B(module_3_W_1_), .Y(_15683_) );
NOR2X1 NOR2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_0_), .B(module_3_W_1_), .Y(_15694_) );
NOR3X1 NOR3X1_471 ( .gnd(gnd), .vdd(vdd), .A(_15672_), .B(_15694_), .C(_15683_), .Y(_15705_) );
OAI21X1 OAI21X1_2586 ( .gnd(gnd), .vdd(vdd), .A(_15705_), .B(_15661_), .C(_15628_), .Y(_15716_) );
INVX1 INVX1_2258 ( .gnd(gnd), .vdd(vdd), .A(_15628_), .Y(_15726_) );
OAI21X1 OAI21X1_2587 ( .gnd(gnd), .vdd(vdd), .A(_15683_), .B(_15694_), .C(_15672_), .Y(_15737_) );
NAND3X1 NAND3X1_3747 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_17_), .B(_15639_), .C(_15650_), .Y(_15748_) );
NAND3X1 NAND3X1_3748 ( .gnd(gnd), .vdd(vdd), .A(_15737_), .B(_15748_), .C(_15726_), .Y(_15759_) );
NAND2X1 NAND2X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_15759_), .B(_15716_), .Y(_15770_) );
NAND2X1 NAND2X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_15606_), .B(_15770_), .Y(_15781_) );
OR2X2 OR2X2_381 ( .gnd(gnd), .vdd(vdd), .A(_15770_), .B(_15606_), .Y(_15792_) );
NAND2X1 NAND2X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_15781_), .B(_15792_), .Y(_15803_) );
XNOR2X1 XNOR2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_15803_), .B(_15595_), .Y(_15814_) );
XNOR2X1 XNOR2X1_430 ( .gnd(gnd), .vdd(vdd), .A(_15814_), .B(bloque_datos[17]), .Y(_15825_) );
AND2X2 AND2X2_359 ( .gnd(gnd), .vdd(vdd), .A(_15825_), .B(_15584_), .Y(_15836_) );
NOR2X1 NOR2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_15584_), .B(_15825_), .Y(_15847_) );
OAI21X1 OAI21X1_2588 ( .gnd(gnd), .vdd(vdd), .A(_15836_), .B(_15847_), .C(_15573_), .Y(_15858_) );
OR2X2 OR2X2_382 ( .gnd(gnd), .vdd(vdd), .A(_15836_), .B(_15847_), .Y(_15869_) );
NOR2X1 NOR2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_15573_), .B(_15869_), .Y(_15880_) );
INVX1 INVX1_2259 ( .gnd(gnd), .vdd(vdd), .A(_15880_), .Y(_15891_) );
NAND2X1 NAND2X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_15858_), .B(_15891_), .Y(_15902_) );
AND2X2 AND2X2_360 ( .gnd(gnd), .vdd(vdd), .A(_15902_), .B(_15562_), .Y(_15913_) );
NOR2X1 NOR2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_15562_), .B(_15902_), .Y(_15924_) );
OAI21X1 OAI21X1_2589 ( .gnd(gnd), .vdd(vdd), .A(_15913_), .B(_15924_), .C(_15551_), .Y(_15935_) );
OR2X2 OR2X2_383 ( .gnd(gnd), .vdd(vdd), .A(_15913_), .B(_15924_), .Y(_15946_) );
NOR2X1 NOR2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_15551_), .B(_15946_), .Y(_15957_) );
INVX1 INVX1_2260 ( .gnd(gnd), .vdd(vdd), .A(_15957_), .Y(_15968_) );
NAND2X1 NAND2X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_15935_), .B(_15968_), .Y(_15979_) );
AND2X2 AND2X2_361 ( .gnd(gnd), .vdd(vdd), .A(_15979_), .B(_15540_), .Y(_15990_) );
NOR2X1 NOR2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_15540_), .B(_15979_), .Y(_16001_) );
NOR2X1 NOR2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_16001_), .B(_15990_), .Y(_16012_) );
XNOR2X1 XNOR2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_16012_), .B(bloque_datos_65_bF_buf0_), .Y(_16023_) );
AND2X2 AND2X2_362 ( .gnd(gnd), .vdd(vdd), .A(_16023_), .B(_15529_), .Y(_16034_) );
NOR2X1 NOR2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_15529_), .B(_16023_), .Y(_16045_) );
NOR2X1 NOR2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_16045_), .B(_16034_), .Y(_16056_) );
NOR2X1 NOR2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf1_), .B(_16056_), .Y(_16066_) );
INVX1 INVX1_2261 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf0_), .Y(_16077_) );
INVX1 INVX1_2262 ( .gnd(gnd), .vdd(vdd), .A(_16056_), .Y(_16088_) );
NOR2X1 NOR2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_16077_), .B(_16088_), .Y(_16099_) );
OAI21X1 OAI21X1_2590 ( .gnd(gnd), .vdd(vdd), .A(_16099_), .B(_16066_), .C(_15518_), .Y(_16110_) );
OR2X2 OR2X2_384 ( .gnd(gnd), .vdd(vdd), .A(_16099_), .B(_16066_), .Y(_16121_) );
NOR2X1 NOR2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_15518_), .B(_16121_), .Y(_16132_) );
INVX2 INVX2_546 ( .gnd(gnd), .vdd(vdd), .A(_16132_), .Y(_16143_) );
NAND2X1 NAND2X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_16143_), .Y(_16154_) );
INVX2 INVX2_547 ( .gnd(gnd), .vdd(vdd), .A(_16154_), .Y(_16165_) );
NOR2X1 NOR2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_129_), .B(_16165_), .Y(_16176_) );
AND2X2 AND2X2_363 ( .gnd(gnd), .vdd(vdd), .A(_16165_), .B(module_3_W_129_), .Y(_16187_) );
OAI21X1 OAI21X1_2591 ( .gnd(gnd), .vdd(vdd), .A(_16187_), .B(_16176_), .C(_15496_), .Y(_16198_) );
OR2X2 OR2X2_385 ( .gnd(gnd), .vdd(vdd), .A(_16187_), .B(_16176_), .Y(_16209_) );
OR2X2 OR2X2_386 ( .gnd(gnd), .vdd(vdd), .A(_16209_), .B(_15496_), .Y(_16220_) );
NAND2X1 NAND2X1_2131 ( .gnd(gnd), .vdd(vdd), .A(_16198_), .B(_16220_), .Y(_16231_) );
NAND2X1 NAND2X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_15474_), .B(_16231_), .Y(_16242_) );
NOR2X1 NOR2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_15474_), .B(_16231_), .Y(_16253_) );
INVX1 INVX1_2263 ( .gnd(gnd), .vdd(vdd), .A(_16253_), .Y(_16264_) );
NAND2X1 NAND2X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_16242_), .B(_16264_), .Y(_16275_) );
NAND2X1 NAND2X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_15463_), .B(_16275_), .Y(_16286_) );
NOR2X1 NOR2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_15463_), .B(_16275_), .Y(_16297_) );
INVX1 INVX1_2264 ( .gnd(gnd), .vdd(vdd), .A(_16297_), .Y(_16308_) );
NAND2X1 NAND2X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_16286_), .B(_16308_), .Y(_16315_) );
NAND2X1 NAND2X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_15441_), .B(_16315_), .Y(_16316_) );
NOR2X1 NOR2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_15441_), .B(_16315_), .Y(_16317_) );
INVX1 INVX1_2265 ( .gnd(gnd), .vdd(vdd), .A(_16317_), .Y(_16318_) );
NAND2X1 NAND2X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_16316_), .B(_16318_), .Y(_16319_) );
NAND2X1 NAND2X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_15430_), .B(_16319_), .Y(_16320_) );
NOR2X1 NOR2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_15430_), .B(_16319_), .Y(_16321_) );
INVX1 INVX1_2266 ( .gnd(gnd), .vdd(vdd), .A(_16321_), .Y(_16322_) );
NAND2X1 NAND2X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_16320_), .B(_16322_), .Y(_16323_) );
INVX2 INVX2_548 ( .gnd(gnd), .vdd(vdd), .A(_16323_), .Y(_16324_) );
NOR2X1 NOR2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_177_), .B(_16324_), .Y(_16325_) );
NAND2X1 NAND2X1_2140 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_177_), .B(_16324_), .Y(_16326_) );
INVX2 INVX2_549 ( .gnd(gnd), .vdd(vdd), .A(_16326_), .Y(_16327_) );
OAI21X1 OAI21X1_2592 ( .gnd(gnd), .vdd(vdd), .A(_16327_), .B(_16325_), .C(_15408_), .Y(_16328_) );
OR2X2 OR2X2_387 ( .gnd(gnd), .vdd(vdd), .A(_16327_), .B(_16325_), .Y(_16329_) );
NOR2X1 NOR2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_15408_), .B(_16329_), .Y(_16330_) );
INVX1 INVX1_2267 ( .gnd(gnd), .vdd(vdd), .A(_16330_), .Y(_16331_) );
NAND2X1 NAND2X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_16328_), .B(_16331_), .Y(_16332_) );
NAND2X1 NAND2X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_15386_), .B(_16332_), .Y(_16333_) );
NOR2X1 NOR2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_15386_), .B(_16332_), .Y(_16334_) );
INVX1 INVX1_2268 ( .gnd(gnd), .vdd(vdd), .A(_16334_), .Y(_16335_) );
NAND2X1 NAND2X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_16333_), .B(_16335_), .Y(_16336_) );
NAND2X1 NAND2X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_15375_), .B(_16336_), .Y(_16337_) );
NOR2X1 NOR2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_15375_), .B(_16336_), .Y(_16338_) );
INVX1 INVX1_2269 ( .gnd(gnd), .vdd(vdd), .A(_16338_), .Y(_16339_) );
NAND2X1 NAND2X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_16337_), .B(_16339_), .Y(_16340_) );
INVX2 INVX2_550 ( .gnd(gnd), .vdd(vdd), .A(_16340_), .Y(_16341_) );
NOR2X1 NOR2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_209_), .B(_16341_), .Y(_16342_) );
NAND2X1 NAND2X1_2146 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_209_), .B(_16341_), .Y(_16343_) );
INVX2 INVX2_551 ( .gnd(gnd), .vdd(vdd), .A(_16343_), .Y(_16344_) );
OAI21X1 OAI21X1_2593 ( .gnd(gnd), .vdd(vdd), .A(_16344_), .B(_16342_), .C(_15354_), .Y(_16345_) );
OR2X2 OR2X2_388 ( .gnd(gnd), .vdd(vdd), .A(_16344_), .B(_16342_), .Y(_16346_) );
NOR2X1 NOR2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_15354_), .B(_16346_), .Y(_16347_) );
INVX2 INVX2_552 ( .gnd(gnd), .vdd(vdd), .A(_16347_), .Y(_16348_) );
NAND2X1 NAND2X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_16345_), .B(_16348_), .Y(_16349_) );
NAND2X1 NAND2X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_15332_), .B(_16349_), .Y(_16350_) );
NOR2X1 NOR2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_15332_), .B(_16349_), .Y(_16351_) );
INVX1 INVX1_2270 ( .gnd(gnd), .vdd(vdd), .A(_16351_), .Y(_16352_) );
NAND2X1 NAND2X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_16350_), .B(_16352_), .Y(_16353_) );
NAND2X1 NAND2X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_15321_), .B(_16353_), .Y(_16354_) );
NOR2X1 NOR2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_15321_), .B(_16353_), .Y(_16355_) );
INVX1 INVX1_2271 ( .gnd(gnd), .vdd(vdd), .A(_16355_), .Y(_16356_) );
NAND2X1 NAND2X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_16354_), .B(_16356_), .Y(_16357_) );
NOR2X1 NOR2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_14864_), .B(_16357_), .Y(_16358_) );
INVX1 INVX1_2272 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_242_), .Y(_16359_) );
INVX1 INVX1_2273 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_194_), .Y(_16360_) );
INVX1 INVX1_2274 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_178_), .Y(_16361_) );
INVX1 INVX1_2275 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_162_), .Y(_16362_) );
NOR2X1 NOR2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_15496_), .B(_16209_), .Y(_16363_) );
AND2X2 AND2X2_364 ( .gnd(gnd), .vdd(vdd), .A(_16012_), .B(bloque_datos_65_bF_buf3_), .Y(_16364_) );
INVX1 INVX1_2276 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf1_), .Y(_16365_) );
INVX1 INVX1_2277 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf1_), .Y(_16366_) );
INVX1 INVX1_2278 ( .gnd(gnd), .vdd(vdd), .A(_15847_), .Y(_16367_) );
NAND2X1 NAND2X1_2152 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .B(_15814_), .Y(_16368_) );
INVX1 INVX1_2279 ( .gnd(gnd), .vdd(vdd), .A(_15595_), .Y(_16369_) );
NOR2X1 NOR2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_16369_), .B(_15803_), .Y(_16370_) );
INVX1 INVX1_2280 ( .gnd(gnd), .vdd(vdd), .A(_15792_), .Y(_16371_) );
INVX1 INVX1_2281 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf3_), .Y(_16372_) );
INVX1 INVX1_2282 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_18_), .Y(_16373_) );
NAND3X1 NAND3X1_3749 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_2_), .B(module_3_W_0_), .C(module_3_W_1_), .Y(_16374_) );
INVX2 INVX2_553 ( .gnd(gnd), .vdd(vdd), .A(_16374_), .Y(_16375_) );
AOI21X1 AOI21X1_2282 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_0_), .B(module_3_W_1_), .C(module_3_W_2_), .Y(_16376_) );
OAI21X1 OAI21X1_2594 ( .gnd(gnd), .vdd(vdd), .A(_16375_), .B(_16376_), .C(_16373_), .Y(_16377_) );
INVX2 INVX2_554 ( .gnd(gnd), .vdd(vdd), .A(_16376_), .Y(_16378_) );
NAND3X1 NAND3X1_3750 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_18_), .B(_16374_), .C(_16378_), .Y(_16379_) );
NAND3X1 NAND3X1_3751 ( .gnd(gnd), .vdd(vdd), .A(_15705_), .B(_16379_), .C(_16377_), .Y(_16380_) );
AOI21X1 AOI21X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_16374_), .B(_16378_), .C(module_3_W_18_), .Y(_16381_) );
NOR3X1 NOR3X1_472 ( .gnd(gnd), .vdd(vdd), .A(_16373_), .B(_16376_), .C(_16375_), .Y(_16382_) );
OAI21X1 OAI21X1_2595 ( .gnd(gnd), .vdd(vdd), .A(_16382_), .B(_16381_), .C(_15748_), .Y(_16383_) );
NAND2X1 NAND2X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_16380_), .B(_16383_), .Y(_16384_) );
NOR2X1 NOR2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_15759_), .B(_16384_), .Y(_16385_) );
INVX1 INVX1_2283 ( .gnd(gnd), .vdd(vdd), .A(_15759_), .Y(_16386_) );
AOI21X1 AOI21X1_2284 ( .gnd(gnd), .vdd(vdd), .A(_16380_), .B(_16383_), .C(_16386_), .Y(_16387_) );
OAI21X1 OAI21X1_2596 ( .gnd(gnd), .vdd(vdd), .A(_16385_), .B(_16387_), .C(_16372_), .Y(_16388_) );
OR2X2 OR2X2_389 ( .gnd(gnd), .vdd(vdd), .A(_16384_), .B(_15759_), .Y(_16389_) );
INVX1 INVX1_2284 ( .gnd(gnd), .vdd(vdd), .A(_16387_), .Y(_16390_) );
NAND3X1 NAND3X1_3752 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf2_), .B(_16390_), .C(_16389_), .Y(_16391_) );
NAND3X1 NAND3X1_3753 ( .gnd(gnd), .vdd(vdd), .A(_16371_), .B(_16388_), .C(_16391_), .Y(_16392_) );
AOI21X1 AOI21X1_2285 ( .gnd(gnd), .vdd(vdd), .A(_16390_), .B(_16389_), .C(bloque_datos_2_bF_buf1_), .Y(_16393_) );
NOR3X1 NOR3X1_473 ( .gnd(gnd), .vdd(vdd), .A(_16372_), .B(_16387_), .C(_16385_), .Y(_16394_) );
OAI21X1 OAI21X1_2597 ( .gnd(gnd), .vdd(vdd), .A(_16393_), .B(_16394_), .C(_15792_), .Y(_16395_) );
NAND3X1 NAND3X1_3754 ( .gnd(gnd), .vdd(vdd), .A(_16370_), .B(_16392_), .C(_16395_), .Y(_16396_) );
AOI21X1 AOI21X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_16392_), .B(_16395_), .C(_16370_), .Y(_16397_) );
INVX1 INVX1_2285 ( .gnd(gnd), .vdd(vdd), .A(_16397_), .Y(_16398_) );
AOI21X1 AOI21X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_16396_), .B(_16398_), .C(bloque_datos[18]), .Y(_16399_) );
INVX1 INVX1_2286 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .Y(_16400_) );
INVX1 INVX1_2287 ( .gnd(gnd), .vdd(vdd), .A(_16370_), .Y(_16401_) );
NOR3X1 NOR3X1_474 ( .gnd(gnd), .vdd(vdd), .A(_16394_), .B(_15792_), .C(_16393_), .Y(_16402_) );
AOI21X1 AOI21X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_16388_), .B(_16391_), .C(_16371_), .Y(_16403_) );
NOR3X1 NOR3X1_475 ( .gnd(gnd), .vdd(vdd), .A(_16401_), .B(_16403_), .C(_16402_), .Y(_16404_) );
NOR3X1 NOR3X1_476 ( .gnd(gnd), .vdd(vdd), .A(_16400_), .B(_16397_), .C(_16404_), .Y(_16405_) );
NOR3X1 NOR3X1_477 ( .gnd(gnd), .vdd(vdd), .A(_16368_), .B(_16405_), .C(_16399_), .Y(_16406_) );
INVX1 INVX1_2288 ( .gnd(gnd), .vdd(vdd), .A(_16368_), .Y(_16407_) );
OAI21X1 OAI21X1_2598 ( .gnd(gnd), .vdd(vdd), .A(_16404_), .B(_16397_), .C(_16400_), .Y(_16408_) );
INVX2 INVX2_555 ( .gnd(gnd), .vdd(vdd), .A(_16405_), .Y(_16409_) );
AOI21X1 AOI21X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_16408_), .B(_16409_), .C(_16407_), .Y(_16410_) );
NOR3X1 NOR3X1_478 ( .gnd(gnd), .vdd(vdd), .A(_16367_), .B(_16406_), .C(_16410_), .Y(_16411_) );
NAND3X1 NAND3X1_3755 ( .gnd(gnd), .vdd(vdd), .A(_16407_), .B(_16408_), .C(_16409_), .Y(_16412_) );
OAI21X1 OAI21X1_2599 ( .gnd(gnd), .vdd(vdd), .A(_16399_), .B(_16405_), .C(_16368_), .Y(_16413_) );
AOI21X1 AOI21X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_16413_), .B(_16412_), .C(_15847_), .Y(_16414_) );
OAI21X1 OAI21X1_2600 ( .gnd(gnd), .vdd(vdd), .A(_16411_), .B(_16414_), .C(_16366_), .Y(_16415_) );
NAND3X1 NAND3X1_3756 ( .gnd(gnd), .vdd(vdd), .A(_15847_), .B(_16413_), .C(_16412_), .Y(_16416_) );
OAI21X1 OAI21X1_2601 ( .gnd(gnd), .vdd(vdd), .A(_16410_), .B(_16406_), .C(_16367_), .Y(_16417_) );
NAND3X1 NAND3X1_3757 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf0_), .B(_16416_), .C(_16417_), .Y(_16418_) );
NAND3X1 NAND3X1_3758 ( .gnd(gnd), .vdd(vdd), .A(_15880_), .B(_16418_), .C(_16415_), .Y(_16419_) );
AOI21X1 AOI21X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_16416_), .B(_16417_), .C(bloque_datos_34_bF_buf4_), .Y(_16420_) );
NOR3X1 NOR3X1_479 ( .gnd(gnd), .vdd(vdd), .A(_16366_), .B(_16414_), .C(_16411_), .Y(_16421_) );
OAI21X1 OAI21X1_2602 ( .gnd(gnd), .vdd(vdd), .A(_16421_), .B(_16420_), .C(_15891_), .Y(_16422_) );
NAND3X1 NAND3X1_3759 ( .gnd(gnd), .vdd(vdd), .A(_15924_), .B(_16419_), .C(_16422_), .Y(_16423_) );
AOI21X1 AOI21X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_16419_), .B(_16422_), .C(_15924_), .Y(_16424_) );
INVX1 INVX1_2289 ( .gnd(gnd), .vdd(vdd), .A(_16424_), .Y(_16425_) );
AOI21X1 AOI21X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_16423_), .B(_16425_), .C(bloque_datos_50_bF_buf0_), .Y(_16426_) );
INVX1 INVX1_2290 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_50_bF_buf3_), .Y(_16427_) );
INVX1 INVX1_2291 ( .gnd(gnd), .vdd(vdd), .A(_16423_), .Y(_16428_) );
NOR3X1 NOR3X1_480 ( .gnd(gnd), .vdd(vdd), .A(_16427_), .B(_16424_), .C(_16428_), .Y(_16429_) );
NOR2X1 NOR2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_16426_), .B(_16429_), .Y(_16430_) );
NAND2X1 NAND2X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_15957_), .B(_16430_), .Y(_16431_) );
OAI21X1 OAI21X1_2603 ( .gnd(gnd), .vdd(vdd), .A(_16429_), .B(_16426_), .C(_15968_), .Y(_16432_) );
NAND3X1 NAND3X1_3760 ( .gnd(gnd), .vdd(vdd), .A(_16001_), .B(_16432_), .C(_16431_), .Y(_16433_) );
INVX2 INVX2_556 ( .gnd(gnd), .vdd(vdd), .A(_16433_), .Y(_16434_) );
AOI21X1 AOI21X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_16432_), .B(_16431_), .C(_16001_), .Y(_16435_) );
OAI21X1 OAI21X1_2604 ( .gnd(gnd), .vdd(vdd), .A(_16434_), .B(_16435_), .C(_16365_), .Y(_16436_) );
INVX1 INVX1_2292 ( .gnd(gnd), .vdd(vdd), .A(_16001_), .Y(_16437_) );
AND2X2 AND2X2_365 ( .gnd(gnd), .vdd(vdd), .A(_16430_), .B(_15957_), .Y(_16438_) );
INVX1 INVX1_2293 ( .gnd(gnd), .vdd(vdd), .A(_16432_), .Y(_16439_) );
OAI21X1 OAI21X1_2605 ( .gnd(gnd), .vdd(vdd), .A(_16438_), .B(_16439_), .C(_16437_), .Y(_16440_) );
NAND3X1 NAND3X1_3761 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf0_), .B(_16433_), .C(_16440_), .Y(_16441_) );
NAND3X1 NAND3X1_3762 ( .gnd(gnd), .vdd(vdd), .A(_16364_), .B(_16441_), .C(_16436_), .Y(_16442_) );
INVX1 INVX1_2294 ( .gnd(gnd), .vdd(vdd), .A(_16364_), .Y(_16443_) );
AOI21X1 AOI21X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_16433_), .B(_16440_), .C(bloque_datos_66_bF_buf4_), .Y(_16444_) );
NOR3X1 NOR3X1_481 ( .gnd(gnd), .vdd(vdd), .A(_16365_), .B(_16435_), .C(_16434_), .Y(_16445_) );
OAI21X1 OAI21X1_2606 ( .gnd(gnd), .vdd(vdd), .A(_16445_), .B(_16444_), .C(_16443_), .Y(_16446_) );
NAND3X1 NAND3X1_3763 ( .gnd(gnd), .vdd(vdd), .A(_16045_), .B(_16442_), .C(_16446_), .Y(_16447_) );
INVX2 INVX2_557 ( .gnd(gnd), .vdd(vdd), .A(_16045_), .Y(_16448_) );
NOR3X1 NOR3X1_482 ( .gnd(gnd), .vdd(vdd), .A(_16443_), .B(_16444_), .C(_16445_), .Y(_16449_) );
AOI21X1 AOI21X1_2296 ( .gnd(gnd), .vdd(vdd), .A(_16441_), .B(_16436_), .C(_16364_), .Y(_16450_) );
OAI21X1 OAI21X1_2607 ( .gnd(gnd), .vdd(vdd), .A(_16449_), .B(_16450_), .C(_16448_), .Y(_16451_) );
AOI21X1 AOI21X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_16447_), .B(_16451_), .C(bloque_datos_82_bF_buf3_), .Y(_16452_) );
INVX1 INVX1_2295 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf2_), .Y(_16453_) );
NOR3X1 NOR3X1_483 ( .gnd(gnd), .vdd(vdd), .A(_16448_), .B(_16450_), .C(_16449_), .Y(_16454_) );
AOI21X1 AOI21X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_16442_), .B(_16446_), .C(_16045_), .Y(_16455_) );
NOR3X1 NOR3X1_484 ( .gnd(gnd), .vdd(vdd), .A(_16453_), .B(_16455_), .C(_16454_), .Y(_16456_) );
NOR2X1 NOR2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_16452_), .B(_16456_), .Y(_16457_) );
NAND2X1 NAND2X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_16099_), .B(_16457_), .Y(_16458_) );
OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_16077_), .B(_16088_), .C(_16456_), .D(_16452_), .Y(_16459_) );
NAND3X1 NAND3X1_3764 ( .gnd(gnd), .vdd(vdd), .A(_16132_), .B(_16459_), .C(_16458_), .Y(_16460_) );
AND2X2 AND2X2_366 ( .gnd(gnd), .vdd(vdd), .A(_16457_), .B(_16099_), .Y(_16461_) );
INVX2 INVX2_558 ( .gnd(gnd), .vdd(vdd), .A(_16459_), .Y(_16462_) );
OAI21X1 OAI21X1_2608 ( .gnd(gnd), .vdd(vdd), .A(_16461_), .B(_16462_), .C(_16143_), .Y(_16463_) );
AOI21X1 AOI21X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_16460_), .B(_16463_), .C(module_3_W_130_), .Y(_16464_) );
INVX1 INVX1_2296 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_130_), .Y(_16465_) );
NOR3X1 NOR3X1_485 ( .gnd(gnd), .vdd(vdd), .A(_16462_), .B(_16143_), .C(_16461_), .Y(_16466_) );
AOI21X1 AOI21X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_16459_), .B(_16458_), .C(_16132_), .Y(_16467_) );
NOR3X1 NOR3X1_486 ( .gnd(gnd), .vdd(vdd), .A(_16465_), .B(_16467_), .C(_16466_), .Y(_16468_) );
NOR2X1 NOR2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_16464_), .B(_16468_), .Y(_16469_) );
NAND2X1 NAND2X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_16187_), .B(_16469_), .Y(_16470_) );
NOR2X1 NOR2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_16187_), .B(_16469_), .Y(_16471_) );
INVX1 INVX1_2297 ( .gnd(gnd), .vdd(vdd), .A(_16471_), .Y(_16472_) );
NAND3X1 NAND3X1_3765 ( .gnd(gnd), .vdd(vdd), .A(_16363_), .B(_16470_), .C(_16472_), .Y(_16473_) );
INVX1 INVX1_2298 ( .gnd(gnd), .vdd(vdd), .A(_16470_), .Y(_16474_) );
OAI21X1 OAI21X1_2609 ( .gnd(gnd), .vdd(vdd), .A(_16474_), .B(_16471_), .C(_16220_), .Y(_16475_) );
AOI21X1 AOI21X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_16475_), .B(_16473_), .C(module_3_W_146_), .Y(_16476_) );
INVX1 INVX1_2299 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_146_), .Y(_16477_) );
NOR3X1 NOR3X1_487 ( .gnd(gnd), .vdd(vdd), .A(_16220_), .B(_16471_), .C(_16474_), .Y(_16478_) );
AOI21X1 AOI21X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_16470_), .B(_16472_), .C(_16363_), .Y(_16479_) );
NOR3X1 NOR3X1_488 ( .gnd(gnd), .vdd(vdd), .A(_16478_), .B(_16477_), .C(_16479_), .Y(_16480_) );
NOR2X1 NOR2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_16476_), .B(_16480_), .Y(_16481_) );
NAND2X1 NAND2X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_16253_), .B(_16481_), .Y(_16482_) );
OAI21X1 OAI21X1_2610 ( .gnd(gnd), .vdd(vdd), .A(_16480_), .B(_16476_), .C(_16264_), .Y(_16483_) );
AND2X2 AND2X2_367 ( .gnd(gnd), .vdd(vdd), .A(_16482_), .B(_16483_), .Y(_16484_) );
NAND2X1 NAND2X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_16297_), .B(_16484_), .Y(_16485_) );
INVX1 INVX1_2300 ( .gnd(gnd), .vdd(vdd), .A(_16485_), .Y(_16486_) );
NOR2X1 NOR2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_16297_), .B(_16484_), .Y(_16487_) );
OAI21X1 OAI21X1_2611 ( .gnd(gnd), .vdd(vdd), .A(_16486_), .B(_16487_), .C(_16362_), .Y(_16488_) );
NOR2X1 NOR2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_16487_), .B(_16486_), .Y(_16489_) );
NAND2X1 NAND2X1_2159 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_162_), .B(_16489_), .Y(_16490_) );
NAND3X1 NAND3X1_3766 ( .gnd(gnd), .vdd(vdd), .A(_16317_), .B(_16488_), .C(_16490_), .Y(_16491_) );
INVX1 INVX1_2301 ( .gnd(gnd), .vdd(vdd), .A(_16488_), .Y(_16492_) );
AND2X2 AND2X2_368 ( .gnd(gnd), .vdd(vdd), .A(_16489_), .B(module_3_W_162_), .Y(_16493_) );
OAI21X1 OAI21X1_2612 ( .gnd(gnd), .vdd(vdd), .A(_16493_), .B(_16492_), .C(_16318_), .Y(_16494_) );
NAND3X1 NAND3X1_3767 ( .gnd(gnd), .vdd(vdd), .A(_16321_), .B(_16491_), .C(_16494_), .Y(_16495_) );
INVX2 INVX2_559 ( .gnd(gnd), .vdd(vdd), .A(_16495_), .Y(_16496_) );
AOI21X1 AOI21X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_16491_), .B(_16494_), .C(_16321_), .Y(_16497_) );
OAI21X1 OAI21X1_2613 ( .gnd(gnd), .vdd(vdd), .A(_16496_), .B(_16497_), .C(_16361_), .Y(_16498_) );
NOR2X1 NOR2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_16497_), .B(_16496_), .Y(_16499_) );
NAND2X1 NAND2X1_2160 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_178_), .B(_16499_), .Y(_16500_) );
NAND3X1 NAND3X1_3768 ( .gnd(gnd), .vdd(vdd), .A(_16327_), .B(_16498_), .C(_16500_), .Y(_16501_) );
INVX1 INVX1_2302 ( .gnd(gnd), .vdd(vdd), .A(_16498_), .Y(_16502_) );
INVX1 INVX1_2303 ( .gnd(gnd), .vdd(vdd), .A(_16500_), .Y(_16503_) );
OAI21X1 OAI21X1_2614 ( .gnd(gnd), .vdd(vdd), .A(_16503_), .B(_16502_), .C(_16326_), .Y(_16504_) );
NAND3X1 NAND3X1_3769 ( .gnd(gnd), .vdd(vdd), .A(_16330_), .B(_16501_), .C(_16504_), .Y(_16505_) );
INVX2 INVX2_560 ( .gnd(gnd), .vdd(vdd), .A(_16505_), .Y(_16506_) );
AOI21X1 AOI21X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_16501_), .B(_16504_), .C(_16330_), .Y(_16507_) );
OAI21X1 OAI21X1_2615 ( .gnd(gnd), .vdd(vdd), .A(_16506_), .B(_16507_), .C(_16360_), .Y(_16508_) );
INVX1 INVX1_2304 ( .gnd(gnd), .vdd(vdd), .A(_16508_), .Y(_16509_) );
NOR3X1 NOR3X1_489 ( .gnd(gnd), .vdd(vdd), .A(_16360_), .B(_16507_), .C(_16506_), .Y(_16510_) );
NOR2X1 NOR2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_16510_), .B(_16509_), .Y(_16511_) );
NAND2X1 NAND2X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_16334_), .B(_16511_), .Y(_16512_) );
OAI21X1 OAI21X1_2616 ( .gnd(gnd), .vdd(vdd), .A(_16509_), .B(_16510_), .C(_16335_), .Y(_16513_) );
NAND3X1 NAND3X1_3770 ( .gnd(gnd), .vdd(vdd), .A(_16338_), .B(_16513_), .C(_16512_), .Y(_16514_) );
INVX2 INVX2_561 ( .gnd(gnd), .vdd(vdd), .A(_16514_), .Y(_16515_) );
AOI21X1 AOI21X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_16513_), .B(_16512_), .C(_16338_), .Y(_16516_) );
NOR2X1 NOR2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_16516_), .B(_16515_), .Y(_16517_) );
NOR2X1 NOR2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_210_), .B(_16517_), .Y(_16518_) );
INVX1 INVX1_2305 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_210_), .Y(_16519_) );
NOR3X1 NOR3X1_490 ( .gnd(gnd), .vdd(vdd), .A(_16519_), .B(_16516_), .C(_16515_), .Y(_16520_) );
NOR2X1 NOR2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_16520_), .B(_16518_), .Y(_16521_) );
NAND2X1 NAND2X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_16344_), .B(_16521_), .Y(_16522_) );
INVX1 INVX1_2306 ( .gnd(gnd), .vdd(vdd), .A(_16522_), .Y(_16523_) );
OAI21X1 OAI21X1_2617 ( .gnd(gnd), .vdd(vdd), .A(_16518_), .B(_16520_), .C(_16343_), .Y(_16524_) );
INVX2 INVX2_562 ( .gnd(gnd), .vdd(vdd), .A(_16524_), .Y(_16525_) );
NOR2X1 NOR2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_16525_), .B(_16523_), .Y(_16526_) );
NAND2X1 NAND2X1_2163 ( .gnd(gnd), .vdd(vdd), .A(_16347_), .B(_16526_), .Y(_16527_) );
OAI21X1 OAI21X1_2618 ( .gnd(gnd), .vdd(vdd), .A(_16523_), .B(_16525_), .C(_16348_), .Y(_16528_) );
AOI21X1 AOI21X1_2306 ( .gnd(gnd), .vdd(vdd), .A(_16528_), .B(_16527_), .C(module_3_W_226_), .Y(_16529_) );
INVX1 INVX1_2307 ( .gnd(gnd), .vdd(vdd), .A(_16529_), .Y(_16530_) );
NAND3X1 NAND3X1_3771 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_226_), .B(_16528_), .C(_16527_), .Y(_16531_) );
NAND3X1 NAND3X1_3772 ( .gnd(gnd), .vdd(vdd), .A(_16351_), .B(_16531_), .C(_16530_), .Y(_16532_) );
INVX2 INVX2_563 ( .gnd(gnd), .vdd(vdd), .A(_16531_), .Y(_16533_) );
OAI21X1 OAI21X1_2619 ( .gnd(gnd), .vdd(vdd), .A(_16533_), .B(_16529_), .C(_16352_), .Y(_16534_) );
NAND3X1 NAND3X1_3773 ( .gnd(gnd), .vdd(vdd), .A(_16355_), .B(_16534_), .C(_16532_), .Y(_16535_) );
INVX1 INVX1_2308 ( .gnd(gnd), .vdd(vdd), .A(_16535_), .Y(_16536_) );
AOI21X1 AOI21X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_16534_), .B(_16532_), .C(_16355_), .Y(_16537_) );
OAI21X1 OAI21X1_2620 ( .gnd(gnd), .vdd(vdd), .A(_16536_), .B(_16537_), .C(_16359_), .Y(_16538_) );
NOR2X1 NOR2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_16537_), .B(_16536_), .Y(_16539_) );
NAND2X1 NAND2X1_2164 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_242_), .B(_16539_), .Y(_16540_) );
NAND3X1 NAND3X1_3774 ( .gnd(gnd), .vdd(vdd), .A(_16358_), .B(_16538_), .C(_16540_), .Y(_16541_) );
NAND2X1 NAND2X1_2165 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_224_), .B(_15299_), .Y(_16542_) );
OR2X2 OR2X2_390 ( .gnd(gnd), .vdd(vdd), .A(_15299_), .B(module_3_W_224_), .Y(_16543_) );
NAND2X1 NAND2X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_16542_), .B(_16543_), .Y(_16544_) );
INVX4 INVX4_14 ( .gnd(gnd), .vdd(vdd), .A(_16544_), .Y(_16545_) );
INVX2 INVX2_564 ( .gnd(gnd), .vdd(vdd), .A(_16357_), .Y(_16546_) );
NOR2X1 NOR2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_241_), .B(_16546_), .Y(_16547_) );
NOR2X1 NOR2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_16358_), .B(_16547_), .Y(_16548_) );
OAI21X1 OAI21X1_2621 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_240_), .B(_16545_), .C(_16548_), .Y(_16549_) );
INVX1 INVX1_2309 ( .gnd(gnd), .vdd(vdd), .A(_16358_), .Y(_16550_) );
INVX1 INVX1_2310 ( .gnd(gnd), .vdd(vdd), .A(_16538_), .Y(_16551_) );
INVX1 INVX1_2311 ( .gnd(gnd), .vdd(vdd), .A(_16540_), .Y(_16552_) );
OAI21X1 OAI21X1_2622 ( .gnd(gnd), .vdd(vdd), .A(_16552_), .B(_16551_), .C(_16550_), .Y(_16553_) );
INVX1 INVX1_2312 ( .gnd(gnd), .vdd(vdd), .A(_16553_), .Y(_16554_) );
OAI21X1 OAI21X1_2623 ( .gnd(gnd), .vdd(vdd), .A(_16554_), .B(_16549_), .C(_16541_), .Y(_16555_) );
INVX1 INVX1_2313 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_243_), .Y(_16556_) );
NAND2X1 NAND2X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_16532_), .B(_16535_), .Y(_16557_) );
INVX1 INVX1_2314 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_227_), .Y(_16558_) );
OAI21X1 OAI21X1_2624 ( .gnd(gnd), .vdd(vdd), .A(_16348_), .B(_16525_), .C(_16522_), .Y(_16559_) );
INVX1 INVX1_2315 ( .gnd(gnd), .vdd(vdd), .A(_16520_), .Y(_16560_) );
INVX1 INVX1_2316 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_211_), .Y(_16561_) );
INVX1 INVX1_2317 ( .gnd(gnd), .vdd(vdd), .A(_16512_), .Y(_16562_) );
AOI21X1 AOI21X1_2308 ( .gnd(gnd), .vdd(vdd), .A(_16338_), .B(_16513_), .C(_16562_), .Y(_16563_) );
INVX1 INVX1_2318 ( .gnd(gnd), .vdd(vdd), .A(_16510_), .Y(_16564_) );
INVX1 INVX1_2319 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_195_), .Y(_16565_) );
AND2X2 AND2X2_369 ( .gnd(gnd), .vdd(vdd), .A(_16505_), .B(_16501_), .Y(_16566_) );
INVX1 INVX1_2320 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_179_), .Y(_16567_) );
INVX1 INVX1_2321 ( .gnd(gnd), .vdd(vdd), .A(_16491_), .Y(_16568_) );
INVX1 INVX1_2322 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_163_), .Y(_16569_) );
INVX1 INVX1_2323 ( .gnd(gnd), .vdd(vdd), .A(_16483_), .Y(_16570_) );
OAI21X1 OAI21X1_2625 ( .gnd(gnd), .vdd(vdd), .A(_16308_), .B(_16570_), .C(_16482_), .Y(_16571_) );
INVX1 INVX1_2324 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_147_), .Y(_16572_) );
OAI21X1 OAI21X1_2626 ( .gnd(gnd), .vdd(vdd), .A(_16220_), .B(_16471_), .C(_16470_), .Y(_16573_) );
INVX1 INVX1_2325 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_131_), .Y(_16574_) );
OAI21X1 OAI21X1_2627 ( .gnd(gnd), .vdd(vdd), .A(_16143_), .B(_16462_), .C(_16458_), .Y(_16575_) );
OAI21X1 OAI21X1_2628 ( .gnd(gnd), .vdd(vdd), .A(_16450_), .B(_16448_), .C(_16442_), .Y(_16576_) );
OAI21X1 OAI21X1_2629 ( .gnd(gnd), .vdd(vdd), .A(_16439_), .B(_16437_), .C(_16431_), .Y(_16577_) );
INVX1 INVX1_2326 ( .gnd(gnd), .vdd(vdd), .A(_16429_), .Y(_16578_) );
AND2X2 AND2X2_370 ( .gnd(gnd), .vdd(vdd), .A(_16423_), .B(_16419_), .Y(_16579_) );
AOI21X1 AOI21X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_16413_), .B(_15847_), .C(_16406_), .Y(_16580_) );
INVX2 INVX2_565 ( .gnd(gnd), .vdd(vdd), .A(_16580_), .Y(_16581_) );
OAI21X1 OAI21X1_2630 ( .gnd(gnd), .vdd(vdd), .A(_16403_), .B(_16401_), .C(_16392_), .Y(_16582_) );
NOR3X1 NOR3X1_491 ( .gnd(gnd), .vdd(vdd), .A(_16381_), .B(_15748_), .C(_16382_), .Y(_16583_) );
AOI21X1 AOI21X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_16386_), .B(_16383_), .C(_16583_), .Y(_16584_) );
INVX1 INVX1_2327 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_19_), .Y(_16585_) );
INVX2 INVX2_566 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_3_), .Y(_16586_) );
NOR2X1 NOR2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_16586_), .B(_16374_), .Y(_16587_) );
AND2X2 AND2X2_371 ( .gnd(gnd), .vdd(vdd), .A(_16374_), .B(_16586_), .Y(_16588_) );
OAI21X1 OAI21X1_2631 ( .gnd(gnd), .vdd(vdd), .A(_16588_), .B(_16587_), .C(_16585_), .Y(_16589_) );
NOR2X1 NOR2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_16587_), .B(_16588_), .Y(_16590_) );
NAND2X1 NAND2X1_2168 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_19_), .B(_16590_), .Y(_16591_) );
AOI21X1 AOI21X1_2311 ( .gnd(gnd), .vdd(vdd), .A(_16589_), .B(_16591_), .C(_16379_), .Y(_16592_) );
INVX1 INVX1_2328 ( .gnd(gnd), .vdd(vdd), .A(_16587_), .Y(_16593_) );
NAND2X1 NAND2X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_16586_), .B(_16374_), .Y(_16594_) );
AOI21X1 AOI21X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_16594_), .B(_16593_), .C(module_3_W_19_), .Y(_16595_) );
NOR3X1 NOR3X1_492 ( .gnd(gnd), .vdd(vdd), .A(_16587_), .B(_16585_), .C(_16588_), .Y(_16596_) );
NOR3X1 NOR3X1_493 ( .gnd(gnd), .vdd(vdd), .A(_16382_), .B(_16596_), .C(_16595_), .Y(_16597_) );
OAI21X1 OAI21X1_2632 ( .gnd(gnd), .vdd(vdd), .A(_16592_), .B(_16597_), .C(_16584_), .Y(_16598_) );
NOR2X1 NOR2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_16597_), .B(_16592_), .Y(_16599_) );
OAI21X1 OAI21X1_2633 ( .gnd(gnd), .vdd(vdd), .A(_16385_), .B(_16583_), .C(_16599_), .Y(_16600_) );
AOI21X1 AOI21X1_2313 ( .gnd(gnd), .vdd(vdd), .A(_16598_), .B(_16600_), .C(bloque_datos_3_bF_buf3_), .Y(_16601_) );
INVX1 INVX1_2329 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf2_), .Y(_16602_) );
INVX1 INVX1_2330 ( .gnd(gnd), .vdd(vdd), .A(_16598_), .Y(_16603_) );
AOI21X1 AOI21X1_2314 ( .gnd(gnd), .vdd(vdd), .A(_16379_), .B(_16377_), .C(_15705_), .Y(_16604_) );
OAI21X1 OAI21X1_2634 ( .gnd(gnd), .vdd(vdd), .A(_16604_), .B(_15759_), .C(_16380_), .Y(_16605_) );
AND2X2 AND2X2_372 ( .gnd(gnd), .vdd(vdd), .A(_16599_), .B(_16605_), .Y(_16606_) );
NOR3X1 NOR3X1_494 ( .gnd(gnd), .vdd(vdd), .A(_16603_), .B(_16602_), .C(_16606_), .Y(_16607_) );
OAI21X1 OAI21X1_2635 ( .gnd(gnd), .vdd(vdd), .A(_16607_), .B(_16601_), .C(_16394_), .Y(_16608_) );
OAI21X1 OAI21X1_2636 ( .gnd(gnd), .vdd(vdd), .A(_16606_), .B(_16603_), .C(_16602_), .Y(_16609_) );
NAND3X1 NAND3X1_3775 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf1_), .B(_16598_), .C(_16600_), .Y(_16610_) );
NAND3X1 NAND3X1_3776 ( .gnd(gnd), .vdd(vdd), .A(_16391_), .B(_16610_), .C(_16609_), .Y(_16611_) );
AOI21X1 AOI21X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_16611_), .B(_16608_), .C(_16582_), .Y(_16612_) );
INVX2 INVX2_567 ( .gnd(gnd), .vdd(vdd), .A(_16612_), .Y(_16613_) );
NAND3X1 NAND3X1_3777 ( .gnd(gnd), .vdd(vdd), .A(_16582_), .B(_16611_), .C(_16608_), .Y(_16614_) );
AOI21X1 AOI21X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_16614_), .B(_16613_), .C(bloque_datos_19_bF_buf3_), .Y(_16615_) );
INVX1 INVX1_2331 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf2_), .Y(_16616_) );
INVX2 INVX2_568 ( .gnd(gnd), .vdd(vdd), .A(_16614_), .Y(_16617_) );
NOR3X1 NOR3X1_495 ( .gnd(gnd), .vdd(vdd), .A(_16616_), .B(_16612_), .C(_16617_), .Y(_16618_) );
OAI21X1 OAI21X1_2637 ( .gnd(gnd), .vdd(vdd), .A(_16618_), .B(_16615_), .C(_16405_), .Y(_16619_) );
OAI21X1 OAI21X1_2638 ( .gnd(gnd), .vdd(vdd), .A(_16617_), .B(_16612_), .C(_16616_), .Y(_16620_) );
NAND3X1 NAND3X1_3778 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf1_), .B(_16614_), .C(_16613_), .Y(_16621_) );
NAND3X1 NAND3X1_3779 ( .gnd(gnd), .vdd(vdd), .A(_16409_), .B(_16620_), .C(_16621_), .Y(_16622_) );
AOI21X1 AOI21X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_16622_), .B(_16619_), .C(_16581_), .Y(_16623_) );
NAND2X1 NAND2X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_16622_), .B(_16619_), .Y(_16624_) );
NOR2X1 NOR2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_16580_), .B(_16624_), .Y(_16625_) );
OAI21X1 OAI21X1_2639 ( .gnd(gnd), .vdd(vdd), .A(_16625_), .B(_16623_), .C(bloque_datos_35_bF_buf1_), .Y(_16626_) );
INVX1 INVX1_2332 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf0_), .Y(_16627_) );
INVX1 INVX1_2333 ( .gnd(gnd), .vdd(vdd), .A(_16619_), .Y(_16628_) );
INVX1 INVX1_2334 ( .gnd(gnd), .vdd(vdd), .A(_16622_), .Y(_16629_) );
OAI21X1 OAI21X1_2640 ( .gnd(gnd), .vdd(vdd), .A(_16628_), .B(_16629_), .C(_16580_), .Y(_16630_) );
NAND3X1 NAND3X1_3780 ( .gnd(gnd), .vdd(vdd), .A(_16622_), .B(_16619_), .C(_16581_), .Y(_16631_) );
NAND3X1 NAND3X1_3781 ( .gnd(gnd), .vdd(vdd), .A(_16627_), .B(_16631_), .C(_16630_), .Y(_16632_) );
NAND3X1 NAND3X1_3782 ( .gnd(gnd), .vdd(vdd), .A(_16421_), .B(_16632_), .C(_16626_), .Y(_16633_) );
OAI21X1 OAI21X1_2641 ( .gnd(gnd), .vdd(vdd), .A(_16625_), .B(_16623_), .C(_16627_), .Y(_16634_) );
NAND3X1 NAND3X1_3783 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf4_), .B(_16631_), .C(_16630_), .Y(_16635_) );
NAND3X1 NAND3X1_3784 ( .gnd(gnd), .vdd(vdd), .A(_16418_), .B(_16635_), .C(_16634_), .Y(_16636_) );
NAND2X1 NAND2X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_16633_), .B(_16636_), .Y(_16637_) );
NAND2X1 NAND2X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_16637_), .B(_16579_), .Y(_16638_) );
OR2X2 OR2X2_391 ( .gnd(gnd), .vdd(vdd), .A(_16579_), .B(_16637_), .Y(_16639_) );
NAND2X1 NAND2X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_16638_), .B(_16639_), .Y(_16640_) );
XNOR2X1 XNOR2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_16640_), .B(bloque_datos_51_bF_buf1_), .Y(_16641_) );
OR2X2 OR2X2_392 ( .gnd(gnd), .vdd(vdd), .A(_16641_), .B(_16578_), .Y(_16642_) );
NOR2X1 NOR2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_16424_), .B(_16428_), .Y(_16643_) );
INVX2 INVX2_569 ( .gnd(gnd), .vdd(vdd), .A(_16643_), .Y(_16644_) );
OAI21X1 OAI21X1_2642 ( .gnd(gnd), .vdd(vdd), .A(_16427_), .B(_16644_), .C(_16641_), .Y(_16645_) );
AOI21X1 AOI21X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_16645_), .B(_16642_), .C(_16577_), .Y(_16646_) );
INVX2 INVX2_570 ( .gnd(gnd), .vdd(vdd), .A(_16577_), .Y(_16647_) );
NOR2X1 NOR2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_16578_), .B(_16641_), .Y(_16648_) );
NAND2X1 NAND2X1_2174 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf0_), .B(_16640_), .Y(_16649_) );
OR2X2 OR2X2_393 ( .gnd(gnd), .vdd(vdd), .A(_16640_), .B(bloque_datos_51_bF_buf4_), .Y(_16650_) );
AOI21X1 AOI21X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_16649_), .B(_16650_), .C(_16429_), .Y(_16651_) );
NOR3X1 NOR3X1_496 ( .gnd(gnd), .vdd(vdd), .A(_16647_), .B(_16651_), .C(_16648_), .Y(_16652_) );
OAI21X1 OAI21X1_2643 ( .gnd(gnd), .vdd(vdd), .A(_16646_), .B(_16652_), .C(bloque_datos_67_bF_buf3_), .Y(_16653_) );
INVX1 INVX1_2335 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf2_), .Y(_16654_) );
NOR2X1 NOR2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_16652_), .B(_16646_), .Y(_16655_) );
NAND2X1 NAND2X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_16654_), .B(_16655_), .Y(_16656_) );
NAND3X1 NAND3X1_3785 ( .gnd(gnd), .vdd(vdd), .A(_16445_), .B(_16653_), .C(_16656_), .Y(_16657_) );
OAI21X1 OAI21X1_2644 ( .gnd(gnd), .vdd(vdd), .A(_16646_), .B(_16652_), .C(_16654_), .Y(_16658_) );
NAND2X1 NAND2X1_2176 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf1_), .B(_16655_), .Y(_16659_) );
NAND3X1 NAND3X1_3786 ( .gnd(gnd), .vdd(vdd), .A(_16441_), .B(_16658_), .C(_16659_), .Y(_16660_) );
AOI21X1 AOI21X1_2320 ( .gnd(gnd), .vdd(vdd), .A(_16660_), .B(_16657_), .C(_16576_), .Y(_16661_) );
NAND3X1 NAND3X1_3787 ( .gnd(gnd), .vdd(vdd), .A(_16576_), .B(_16660_), .C(_16657_), .Y(_16662_) );
INVX2 INVX2_571 ( .gnd(gnd), .vdd(vdd), .A(_16662_), .Y(_16663_) );
OAI21X1 OAI21X1_2645 ( .gnd(gnd), .vdd(vdd), .A(_16663_), .B(_16661_), .C(bloque_datos_83_bF_buf5_), .Y(_16664_) );
INVX1 INVX1_2336 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf4_), .Y(_16665_) );
INVX2 INVX2_572 ( .gnd(gnd), .vdd(vdd), .A(_16661_), .Y(_16666_) );
NAND3X1 NAND3X1_3788 ( .gnd(gnd), .vdd(vdd), .A(_16665_), .B(_16662_), .C(_16666_), .Y(_16667_) );
NAND3X1 NAND3X1_3789 ( .gnd(gnd), .vdd(vdd), .A(_16456_), .B(_16667_), .C(_16664_), .Y(_16668_) );
INVX1 INVX1_2337 ( .gnd(gnd), .vdd(vdd), .A(_16456_), .Y(_16669_) );
OAI21X1 OAI21X1_2646 ( .gnd(gnd), .vdd(vdd), .A(_16663_), .B(_16661_), .C(_16665_), .Y(_16670_) );
NAND3X1 NAND3X1_3790 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf3_), .B(_16662_), .C(_16666_), .Y(_16671_) );
NAND3X1 NAND3X1_3791 ( .gnd(gnd), .vdd(vdd), .A(_16669_), .B(_16671_), .C(_16670_), .Y(_16672_) );
AOI21X1 AOI21X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_16668_), .B(_16672_), .C(_16575_), .Y(_16673_) );
NAND3X1 NAND3X1_3792 ( .gnd(gnd), .vdd(vdd), .A(_16575_), .B(_16668_), .C(_16672_), .Y(_16674_) );
INVX2 INVX2_573 ( .gnd(gnd), .vdd(vdd), .A(_16674_), .Y(_16675_) );
OAI21X1 OAI21X1_2647 ( .gnd(gnd), .vdd(vdd), .A(_16675_), .B(_16673_), .C(_16574_), .Y(_16676_) );
INVX1 INVX1_2338 ( .gnd(gnd), .vdd(vdd), .A(_16673_), .Y(_16677_) );
NAND3X1 NAND3X1_3793 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_131_), .B(_16674_), .C(_16677_), .Y(_16678_) );
NAND2X1 NAND2X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_16678_), .B(_16676_), .Y(_16679_) );
NAND2X1 NAND2X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_16468_), .B(_16679_), .Y(_16680_) );
INVX1 INVX1_2339 ( .gnd(gnd), .vdd(vdd), .A(_16468_), .Y(_16681_) );
NAND3X1 NAND3X1_3794 ( .gnd(gnd), .vdd(vdd), .A(_16681_), .B(_16678_), .C(_16676_), .Y(_16682_) );
NAND3X1 NAND3X1_3795 ( .gnd(gnd), .vdd(vdd), .A(_16682_), .B(_16680_), .C(_16573_), .Y(_16683_) );
INVX1 INVX1_2340 ( .gnd(gnd), .vdd(vdd), .A(_16683_), .Y(_16684_) );
AND2X2 AND2X2_373 ( .gnd(gnd), .vdd(vdd), .A(_16680_), .B(_16682_), .Y(_16685_) );
NOR2X1 NOR2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_16573_), .B(_16685_), .Y(_16686_) );
OAI21X1 OAI21X1_2648 ( .gnd(gnd), .vdd(vdd), .A(_16686_), .B(_16684_), .C(_16572_), .Y(_16687_) );
NOR3X1 NOR3X1_497 ( .gnd(gnd), .vdd(vdd), .A(_16572_), .B(_16684_), .C(_16686_), .Y(_16688_) );
INVX2 INVX2_574 ( .gnd(gnd), .vdd(vdd), .A(_16688_), .Y(_16689_) );
NAND3X1 NAND3X1_3796 ( .gnd(gnd), .vdd(vdd), .A(_16480_), .B(_16687_), .C(_16689_), .Y(_16690_) );
INVX1 INVX1_2341 ( .gnd(gnd), .vdd(vdd), .A(_16480_), .Y(_16691_) );
INVX1 INVX1_2342 ( .gnd(gnd), .vdd(vdd), .A(_16687_), .Y(_16692_) );
OAI21X1 OAI21X1_2649 ( .gnd(gnd), .vdd(vdd), .A(_16692_), .B(_16688_), .C(_16691_), .Y(_16693_) );
NAND3X1 NAND3X1_3797 ( .gnd(gnd), .vdd(vdd), .A(_16693_), .B(_16571_), .C(_16690_), .Y(_16694_) );
INVX1 INVX1_2343 ( .gnd(gnd), .vdd(vdd), .A(_16694_), .Y(_16695_) );
AOI21X1 AOI21X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_16693_), .B(_16690_), .C(_16571_), .Y(_16696_) );
OAI21X1 OAI21X1_2650 ( .gnd(gnd), .vdd(vdd), .A(_16695_), .B(_16696_), .C(_16569_), .Y(_16697_) );
NOR2X1 NOR2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_16696_), .B(_16695_), .Y(_16698_) );
NAND2X1 NAND2X1_2179 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_163_), .B(_16698_), .Y(_16699_) );
NAND2X1 NAND2X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_16697_), .B(_16699_), .Y(_16700_) );
NOR2X1 NOR2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_16490_), .B(_16700_), .Y(_16701_) );
INVX2 INVX2_575 ( .gnd(gnd), .vdd(vdd), .A(_16489_), .Y(_16702_) );
OAI21X1 OAI21X1_2651 ( .gnd(gnd), .vdd(vdd), .A(_16362_), .B(_16702_), .C(_16700_), .Y(_16703_) );
INVX2 INVX2_576 ( .gnd(gnd), .vdd(vdd), .A(_16703_), .Y(_16704_) );
NOR2X1 NOR2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_16701_), .B(_16704_), .Y(_16705_) );
OAI21X1 OAI21X1_2652 ( .gnd(gnd), .vdd(vdd), .A(_16496_), .B(_16568_), .C(_16705_), .Y(_16706_) );
AOI21X1 AOI21X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_16321_), .B(_16494_), .C(_16568_), .Y(_16707_) );
OAI21X1 OAI21X1_2653 ( .gnd(gnd), .vdd(vdd), .A(_16704_), .B(_16701_), .C(_16707_), .Y(_16708_) );
NAND2X1 NAND2X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_16708_), .B(_16706_), .Y(_16709_) );
NAND2X1 NAND2X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_16567_), .B(_16709_), .Y(_16710_) );
NOR2X1 NOR2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_16567_), .B(_16709_), .Y(_16711_) );
INVX2 INVX2_577 ( .gnd(gnd), .vdd(vdd), .A(_16711_), .Y(_16712_) );
NAND3X1 NAND3X1_3798 ( .gnd(gnd), .vdd(vdd), .A(_16503_), .B(_16710_), .C(_16712_), .Y(_16713_) );
INVX1 INVX1_2344 ( .gnd(gnd), .vdd(vdd), .A(_16710_), .Y(_16714_) );
OAI21X1 OAI21X1_2654 ( .gnd(gnd), .vdd(vdd), .A(_16714_), .B(_16711_), .C(_16500_), .Y(_16715_) );
NAND2X1 NAND2X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_16715_), .B(_16713_), .Y(_16716_) );
NOR2X1 NOR2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_16566_), .B(_16716_), .Y(_16717_) );
INVX1 INVX1_2345 ( .gnd(gnd), .vdd(vdd), .A(_16713_), .Y(_16718_) );
INVX1 INVX1_2346 ( .gnd(gnd), .vdd(vdd), .A(_16715_), .Y(_16719_) );
OAI21X1 OAI21X1_2655 ( .gnd(gnd), .vdd(vdd), .A(_16718_), .B(_16719_), .C(_16566_), .Y(_16720_) );
INVX1 INVX1_2347 ( .gnd(gnd), .vdd(vdd), .A(_16720_), .Y(_16721_) );
OAI21X1 OAI21X1_2656 ( .gnd(gnd), .vdd(vdd), .A(_16721_), .B(_16717_), .C(_16565_), .Y(_16722_) );
NOR2X1 NOR2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_16717_), .B(_16721_), .Y(_16723_) );
NAND2X1 NAND2X1_2184 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_195_), .B(_16723_), .Y(_16724_) );
NAND2X1 NAND2X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_16722_), .B(_16724_), .Y(_16725_) );
OR2X2 OR2X2_394 ( .gnd(gnd), .vdd(vdd), .A(_16725_), .B(_16564_), .Y(_16726_) );
AOI21X1 AOI21X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_16722_), .B(_16724_), .C(_16510_), .Y(_16727_) );
INVX1 INVX1_2348 ( .gnd(gnd), .vdd(vdd), .A(_16727_), .Y(_16728_) );
NAND2X1 NAND2X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_16728_), .B(_16726_), .Y(_16729_) );
NOR2X1 NOR2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_16563_), .B(_16729_), .Y(_16730_) );
NOR2X1 NOR2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_16564_), .B(_16725_), .Y(_16731_) );
OAI21X1 OAI21X1_2657 ( .gnd(gnd), .vdd(vdd), .A(_16731_), .B(_16727_), .C(_16563_), .Y(_16732_) );
INVX2 INVX2_578 ( .gnd(gnd), .vdd(vdd), .A(_16732_), .Y(_16733_) );
OAI21X1 OAI21X1_2658 ( .gnd(gnd), .vdd(vdd), .A(_16730_), .B(_16733_), .C(_16561_), .Y(_16734_) );
INVX1 INVX1_2349 ( .gnd(gnd), .vdd(vdd), .A(_16734_), .Y(_16735_) );
NOR2X1 NOR2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_16727_), .B(_16731_), .Y(_16736_) );
OAI21X1 OAI21X1_2659 ( .gnd(gnd), .vdd(vdd), .A(_16562_), .B(_16515_), .C(_16736_), .Y(_16737_) );
NAND2X1 NAND2X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_16732_), .B(_16737_), .Y(_16738_) );
NOR2X1 NOR2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_16561_), .B(_16738_), .Y(_16739_) );
NOR3X1 NOR3X1_498 ( .gnd(gnd), .vdd(vdd), .A(_16560_), .B(_16739_), .C(_16735_), .Y(_16740_) );
NOR2X1 NOR2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_16733_), .B(_16730_), .Y(_16741_) );
NAND2X1 NAND2X1_2188 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_211_), .B(_16741_), .Y(_16742_) );
AOI21X1 AOI21X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_16734_), .B(_16742_), .C(_16520_), .Y(_16743_) );
NOR2X1 NOR2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_16743_), .B(_16740_), .Y(_16744_) );
AND2X2 AND2X2_374 ( .gnd(gnd), .vdd(vdd), .A(_16744_), .B(_16559_), .Y(_16745_) );
INVX1 INVX1_2350 ( .gnd(gnd), .vdd(vdd), .A(_16559_), .Y(_16746_) );
OAI21X1 OAI21X1_2660 ( .gnd(gnd), .vdd(vdd), .A(_16740_), .B(_16743_), .C(_16746_), .Y(_16747_) );
INVX2 INVX2_579 ( .gnd(gnd), .vdd(vdd), .A(_16747_), .Y(_16748_) );
OAI21X1 OAI21X1_2661 ( .gnd(gnd), .vdd(vdd), .A(_16745_), .B(_16748_), .C(_16558_), .Y(_16749_) );
NOR2X1 NOR2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_16748_), .B(_16745_), .Y(_16750_) );
NAND2X1 NAND2X1_2189 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_227_), .B(_16750_), .Y(_16751_) );
NAND3X1 NAND3X1_3799 ( .gnd(gnd), .vdd(vdd), .A(_16533_), .B(_16749_), .C(_16751_), .Y(_16752_) );
NAND2X1 NAND2X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_16749_), .B(_16751_), .Y(_16753_) );
NAND2X1 NAND2X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_16531_), .B(_16753_), .Y(_16754_) );
NAND3X1 NAND3X1_3800 ( .gnd(gnd), .vdd(vdd), .A(_16557_), .B(_16752_), .C(_16754_), .Y(_16755_) );
INVX2 INVX2_580 ( .gnd(gnd), .vdd(vdd), .A(_16755_), .Y(_16756_) );
AND2X2 AND2X2_375 ( .gnd(gnd), .vdd(vdd), .A(_16535_), .B(_16532_), .Y(_16757_) );
INVX1 INVX1_2351 ( .gnd(gnd), .vdd(vdd), .A(_16752_), .Y(_16758_) );
AOI21X1 AOI21X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_16749_), .B(_16751_), .C(_16533_), .Y(_16759_) );
OAI21X1 OAI21X1_2662 ( .gnd(gnd), .vdd(vdd), .A(_16758_), .B(_16759_), .C(_16757_), .Y(_16760_) );
INVX2 INVX2_581 ( .gnd(gnd), .vdd(vdd), .A(_16760_), .Y(_16761_) );
OAI21X1 OAI21X1_2663 ( .gnd(gnd), .vdd(vdd), .A(_16761_), .B(_16756_), .C(_16556_), .Y(_16762_) );
NOR2X1 NOR2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_16756_), .B(_16761_), .Y(_16763_) );
NAND2X1 NAND2X1_2192 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_243_), .B(_16763_), .Y(_16764_) );
NAND2X1 NAND2X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_16762_), .B(_16764_), .Y(_16765_) );
OR2X2 OR2X2_395 ( .gnd(gnd), .vdd(vdd), .A(_16765_), .B(_16540_), .Y(_16766_) );
INVX2 INVX2_582 ( .gnd(gnd), .vdd(vdd), .A(_16539_), .Y(_16767_) );
OAI21X1 OAI21X1_2664 ( .gnd(gnd), .vdd(vdd), .A(_16767_), .B(_16359_), .C(_16765_), .Y(_16768_) );
AOI21X1 AOI21X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_16768_), .B(_16766_), .C(_16555_), .Y(_16769_) );
INVX1 INVX1_2352 ( .gnd(gnd), .vdd(vdd), .A(_16555_), .Y(_16770_) );
NAND2X1 NAND2X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_16768_), .B(_16766_), .Y(_16771_) );
NOR2X1 NOR2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_16770_), .B(_16771_), .Y(_16772_) );
NOR2X1 NOR2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_16769_), .B(_16772_), .Y(_16773_) );
INVX2 INVX2_583 ( .gnd(gnd), .vdd(vdd), .A(_16773_), .Y(module_3_H_15_) );
NOR2X1 NOR2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_240_), .B(_16545_), .Y(_16774_) );
OAI21X1 OAI21X1_2665 ( .gnd(gnd), .vdd(vdd), .A(_16547_), .B(_16358_), .C(_16774_), .Y(_16775_) );
NAND2X1 NAND2X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_16775_), .B(_16549_), .Y(_16776_) );
INVX2 INVX2_584 ( .gnd(gnd), .vdd(vdd), .A(_16776_), .Y(module_3_H_13_) );
NAND2X1 NAND2X1_2196 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_240_), .B(_16545_), .Y(_16777_) );
INVX1 INVX1_2353 ( .gnd(gnd), .vdd(vdd), .A(_16777_), .Y(_16778_) );
NOR2X1 NOR2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_16774_), .B(_16778_), .Y(module_3_H_0_) );
INVX1 INVX1_2354 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_0_), .Y(module_3_H_12_) );
INVX1 INVX1_2355 ( .gnd(gnd), .vdd(vdd), .A(_16549_), .Y(_16779_) );
OAI21X1 OAI21X1_2666 ( .gnd(gnd), .vdd(vdd), .A(_16774_), .B(_16778_), .C(module_3_H_13_), .Y(_16780_) );
INVX2 INVX2_585 ( .gnd(gnd), .vdd(vdd), .A(_16780_), .Y(_16781_) );
AOI21X1 AOI21X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_16779_), .B(_16777_), .C(_16781_), .Y(module_3_H_1_) );
NAND3X1 NAND3X1_3801 ( .gnd(gnd), .vdd(vdd), .A(_16541_), .B(_16779_), .C(_16553_), .Y(_16782_) );
INVX1 INVX1_2356 ( .gnd(gnd), .vdd(vdd), .A(_16541_), .Y(_16783_) );
OAI21X1 OAI21X1_2667 ( .gnd(gnd), .vdd(vdd), .A(_16554_), .B(_16783_), .C(_16549_), .Y(_16784_) );
AND2X2 AND2X2_376 ( .gnd(gnd), .vdd(vdd), .A(_16784_), .B(_16782_), .Y(module_3_H_14_) );
NAND2X1 NAND2X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_16781_), .B(module_3_H_14_), .Y(_16785_) );
INVX1 INVX1_2357 ( .gnd(gnd), .vdd(vdd), .A(_16785_), .Y(_16786_) );
NOR2X1 NOR2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_16781_), .B(module_3_H_14_), .Y(_16787_) );
NOR2X1 NOR2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_16787_), .B(_16786_), .Y(module_3_H_2_) );
NOR3X1 NOR3X1_499 ( .gnd(gnd), .vdd(vdd), .A(_16785_), .B(_16769_), .C(_16772_), .Y(_16788_) );
NOR2X1 NOR2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_16786_), .B(_16773_), .Y(_16789_) );
NOR2X1 NOR2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_16788_), .B(_16789_), .Y(module_3_H_3_) );
AOI21X1 AOI21X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_16762_), .B(_16764_), .C(_16552_), .Y(_16790_) );
OAI21X1 OAI21X1_2668 ( .gnd(gnd), .vdd(vdd), .A(_16770_), .B(_16790_), .C(_16766_), .Y(_16791_) );
INVX1 INVX1_2358 ( .gnd(gnd), .vdd(vdd), .A(_16764_), .Y(_16792_) );
AOI21X1 AOI21X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_16557_), .B(_16754_), .C(_16758_), .Y(_16793_) );
OAI21X1 OAI21X1_2669 ( .gnd(gnd), .vdd(vdd), .A(_16735_), .B(_16739_), .C(_16560_), .Y(_16794_) );
AOI21X1 AOI21X1_2331 ( .gnd(gnd), .vdd(vdd), .A(_16559_), .B(_16794_), .C(_16740_), .Y(_16795_) );
INVX1 INVX1_2359 ( .gnd(gnd), .vdd(vdd), .A(_16563_), .Y(_16796_) );
AOI21X1 AOI21X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_16796_), .B(_16728_), .C(_16731_), .Y(_16797_) );
NAND2X1 NAND2X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_16501_), .B(_16505_), .Y(_16798_) );
AOI21X1 AOI21X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_16798_), .B(_16715_), .C(_16718_), .Y(_16799_) );
INVX1 INVX1_2360 ( .gnd(gnd), .vdd(vdd), .A(_16701_), .Y(_16800_) );
OAI21X1 OAI21X1_2670 ( .gnd(gnd), .vdd(vdd), .A(_16704_), .B(_16707_), .C(_16800_), .Y(_16801_) );
INVX1 INVX1_2361 ( .gnd(gnd), .vdd(vdd), .A(_16801_), .Y(_16802_) );
AND2X2 AND2X2_377 ( .gnd(gnd), .vdd(vdd), .A(_16694_), .B(_16690_), .Y(_16803_) );
NAND2X1 NAND2X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_16680_), .B(_16683_), .Y(_16804_) );
AND2X2 AND2X2_378 ( .gnd(gnd), .vdd(vdd), .A(_16674_), .B(_16668_), .Y(_16805_) );
INVX2 INVX2_586 ( .gnd(gnd), .vdd(vdd), .A(_16670_), .Y(_16806_) );
AOI21X1 AOI21X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_16658_), .B(_16659_), .C(_16441_), .Y(_16807_) );
AOI21X1 AOI21X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_16576_), .B(_16660_), .C(_16807_), .Y(_16808_) );
INVX2 INVX2_587 ( .gnd(gnd), .vdd(vdd), .A(_16658_), .Y(_16809_) );
AOI21X1 AOI21X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_16577_), .B(_16645_), .C(_16648_), .Y(_16810_) );
INVX1 INVX1_2362 ( .gnd(gnd), .vdd(vdd), .A(_16640_), .Y(_16811_) );
NOR2X1 NOR2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf3_), .B(_16811_), .Y(_16812_) );
NAND2X1 NAND2X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_16419_), .B(_16423_), .Y(_16813_) );
INVX1 INVX1_2363 ( .gnd(gnd), .vdd(vdd), .A(_16633_), .Y(_16814_) );
AOI21X1 AOI21X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_16636_), .B(_16813_), .C(_16814_), .Y(_16815_) );
INVX2 INVX2_588 ( .gnd(gnd), .vdd(vdd), .A(_16634_), .Y(_16816_) );
AOI21X1 AOI21X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_16622_), .B(_16581_), .C(_16628_), .Y(_16817_) );
AOI21X1 AOI21X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_16610_), .B(_16609_), .C(_16391_), .Y(_16818_) );
AOI21X1 AOI21X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_16611_), .B(_16582_), .C(_16818_), .Y(_16819_) );
OAI21X1 OAI21X1_2671 ( .gnd(gnd), .vdd(vdd), .A(_16595_), .B(_16596_), .C(_16382_), .Y(_16820_) );
OAI21X1 OAI21X1_2672 ( .gnd(gnd), .vdd(vdd), .A(_16584_), .B(_16597_), .C(_16820_), .Y(_16821_) );
INVX1 INVX1_2364 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_4_), .Y(_16822_) );
OAI21X1 OAI21X1_2673 ( .gnd(gnd), .vdd(vdd), .A(_16374_), .B(_16586_), .C(_16822_), .Y(_16823_) );
NAND2X1 NAND2X1_2201 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_4_), .B(_16587_), .Y(_16824_) );
AOI21X1 AOI21X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_16823_), .B(_16824_), .C(_15617_), .Y(_16825_) );
INVX1 INVX1_2365 ( .gnd(gnd), .vdd(vdd), .A(_16823_), .Y(_16826_) );
NOR3X1 NOR3X1_500 ( .gnd(gnd), .vdd(vdd), .A(_16586_), .B(_16822_), .C(_16374_), .Y(_16827_) );
NOR3X1 NOR3X1_501 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_0_), .B(_16827_), .C(_16826_), .Y(_16828_) );
OAI21X1 OAI21X1_2674 ( .gnd(gnd), .vdd(vdd), .A(_16828_), .B(_16825_), .C(module_3_W_20_), .Y(_16829_) );
INVX1 INVX1_2366 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_20_), .Y(_16830_) );
OAI21X1 OAI21X1_2675 ( .gnd(gnd), .vdd(vdd), .A(_16826_), .B(_16827_), .C(module_3_W_0_), .Y(_16831_) );
NAND3X1 NAND3X1_3802 ( .gnd(gnd), .vdd(vdd), .A(_15617_), .B(_16823_), .C(_16824_), .Y(_16832_) );
NAND3X1 NAND3X1_3803 ( .gnd(gnd), .vdd(vdd), .A(_16830_), .B(_16832_), .C(_16831_), .Y(_16833_) );
NAND3X1 NAND3X1_3804 ( .gnd(gnd), .vdd(vdd), .A(_16589_), .B(_16833_), .C(_16829_), .Y(_16834_) );
OAI21X1 OAI21X1_2676 ( .gnd(gnd), .vdd(vdd), .A(_16828_), .B(_16825_), .C(_16830_), .Y(_16835_) );
NAND3X1 NAND3X1_3805 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_20_), .B(_16832_), .C(_16831_), .Y(_16836_) );
NAND3X1 NAND3X1_3806 ( .gnd(gnd), .vdd(vdd), .A(_16595_), .B(_16836_), .C(_16835_), .Y(_16837_) );
NAND3X1 NAND3X1_3807 ( .gnd(gnd), .vdd(vdd), .A(_16834_), .B(_16837_), .C(_16821_), .Y(_16838_) );
NAND3X1 NAND3X1_3808 ( .gnd(gnd), .vdd(vdd), .A(_16379_), .B(_16589_), .C(_16591_), .Y(_16839_) );
AOI21X1 AOI21X1_2342 ( .gnd(gnd), .vdd(vdd), .A(_16839_), .B(_16605_), .C(_16592_), .Y(_16840_) );
NAND3X1 NAND3X1_3809 ( .gnd(gnd), .vdd(vdd), .A(_16595_), .B(_16833_), .C(_16829_), .Y(_16841_) );
NAND3X1 NAND3X1_3810 ( .gnd(gnd), .vdd(vdd), .A(_16589_), .B(_16836_), .C(_16835_), .Y(_16842_) );
NAND3X1 NAND3X1_3811 ( .gnd(gnd), .vdd(vdd), .A(_16840_), .B(_16841_), .C(_16842_), .Y(_16843_) );
XNOR2X1 XNOR2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_14919_), .B(module_3_W_8_), .Y(_16844_) );
INVX1 INVX1_2367 ( .gnd(gnd), .vdd(vdd), .A(_16844_), .Y(_16845_) );
NAND3X1 NAND3X1_3812 ( .gnd(gnd), .vdd(vdd), .A(_16845_), .B(_16843_), .C(_16838_), .Y(_16846_) );
AOI21X1 AOI21X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_16841_), .B(_16842_), .C(_16840_), .Y(_16847_) );
AOI21X1 AOI21X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_16834_), .B(_16837_), .C(_16821_), .Y(_16848_) );
OAI21X1 OAI21X1_2677 ( .gnd(gnd), .vdd(vdd), .A(_16847_), .B(_16848_), .C(_16844_), .Y(_16849_) );
AOI21X1 AOI21X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_16846_), .B(_16849_), .C(bloque_datos_4_bF_buf3_), .Y(_16850_) );
INVX1 INVX1_2368 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf2_), .Y(_16851_) );
NAND3X1 NAND3X1_3813 ( .gnd(gnd), .vdd(vdd), .A(_16844_), .B(_16843_), .C(_16838_), .Y(_16852_) );
OAI21X1 OAI21X1_2678 ( .gnd(gnd), .vdd(vdd), .A(_16847_), .B(_16848_), .C(_16845_), .Y(_16853_) );
AOI21X1 AOI21X1_2346 ( .gnd(gnd), .vdd(vdd), .A(_16852_), .B(_16853_), .C(_16851_), .Y(_16854_) );
OAI21X1 OAI21X1_2679 ( .gnd(gnd), .vdd(vdd), .A(_16850_), .B(_16854_), .C(_16601_), .Y(_16855_) );
NAND3X1 NAND3X1_3814 ( .gnd(gnd), .vdd(vdd), .A(_16851_), .B(_16852_), .C(_16853_), .Y(_16856_) );
NAND3X1 NAND3X1_3815 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf1_), .B(_16846_), .C(_16849_), .Y(_16857_) );
NAND3X1 NAND3X1_3816 ( .gnd(gnd), .vdd(vdd), .A(_16609_), .B(_16856_), .C(_16857_), .Y(_16858_) );
NAND3X1 NAND3X1_3817 ( .gnd(gnd), .vdd(vdd), .A(_16819_), .B(_16858_), .C(_16855_), .Y(_16859_) );
AOI21X1 AOI21X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_16395_), .B(_16370_), .C(_16402_), .Y(_16860_) );
NOR3X1 NOR3X1_502 ( .gnd(gnd), .vdd(vdd), .A(_16394_), .B(_16601_), .C(_16607_), .Y(_16861_) );
OAI21X1 OAI21X1_2680 ( .gnd(gnd), .vdd(vdd), .A(_16861_), .B(_16860_), .C(_16608_), .Y(_16862_) );
OAI21X1 OAI21X1_2681 ( .gnd(gnd), .vdd(vdd), .A(_16850_), .B(_16854_), .C(_16609_), .Y(_16863_) );
NAND3X1 NAND3X1_3818 ( .gnd(gnd), .vdd(vdd), .A(_16601_), .B(_16856_), .C(_16857_), .Y(_16864_) );
NAND3X1 NAND3X1_3819 ( .gnd(gnd), .vdd(vdd), .A(_16864_), .B(_16863_), .C(_16862_), .Y(_16865_) );
NOR2X1 NOR2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_24_), .B(module_3_W_8_), .Y(_16866_) );
INVX1 INVX1_2369 ( .gnd(gnd), .vdd(vdd), .A(_16866_), .Y(_16867_) );
NAND2X1 NAND2X1_2202 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_24_), .B(module_3_W_8_), .Y(_16868_) );
NAND2X1 NAND2X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_16868_), .B(_16867_), .Y(_16869_) );
XNOR2X1 XNOR2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_14941_), .B(_16869_), .Y(_16870_) );
NAND3X1 NAND3X1_3820 ( .gnd(gnd), .vdd(vdd), .A(_16870_), .B(_16859_), .C(_16865_), .Y(_16871_) );
AOI21X1 AOI21X1_2348 ( .gnd(gnd), .vdd(vdd), .A(_16864_), .B(_16863_), .C(_16862_), .Y(_16872_) );
AOI21X1 AOI21X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_16858_), .B(_16855_), .C(_16819_), .Y(_16873_) );
INVX1 INVX1_2370 ( .gnd(gnd), .vdd(vdd), .A(_16870_), .Y(_16874_) );
OAI21X1 OAI21X1_2682 ( .gnd(gnd), .vdd(vdd), .A(_16872_), .B(_16873_), .C(_16874_), .Y(_16875_) );
AOI21X1 AOI21X1_2350 ( .gnd(gnd), .vdd(vdd), .A(_16871_), .B(_16875_), .C(bloque_datos_20_bF_buf3_), .Y(_16876_) );
INVX1 INVX1_2371 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf2_), .Y(_16877_) );
OAI21X1 OAI21X1_2683 ( .gnd(gnd), .vdd(vdd), .A(_16872_), .B(_16873_), .C(_16870_), .Y(_16878_) );
NAND3X1 NAND3X1_3821 ( .gnd(gnd), .vdd(vdd), .A(_16874_), .B(_16859_), .C(_16865_), .Y(_16879_) );
AOI21X1 AOI21X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_16879_), .B(_16878_), .C(_16877_), .Y(_16880_) );
OAI21X1 OAI21X1_2684 ( .gnd(gnd), .vdd(vdd), .A(_16876_), .B(_16880_), .C(_16615_), .Y(_16881_) );
NAND3X1 NAND3X1_3822 ( .gnd(gnd), .vdd(vdd), .A(_16877_), .B(_16879_), .C(_16878_), .Y(_16882_) );
NAND3X1 NAND3X1_3823 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf1_), .B(_16871_), .C(_16875_), .Y(_16883_) );
NAND3X1 NAND3X1_3824 ( .gnd(gnd), .vdd(vdd), .A(_16620_), .B(_16882_), .C(_16883_), .Y(_16884_) );
NAND3X1 NAND3X1_3825 ( .gnd(gnd), .vdd(vdd), .A(_16884_), .B(_16881_), .C(_16817_), .Y(_16885_) );
OAI21X1 OAI21X1_2685 ( .gnd(gnd), .vdd(vdd), .A(_16629_), .B(_16580_), .C(_16619_), .Y(_16886_) );
OAI21X1 OAI21X1_2686 ( .gnd(gnd), .vdd(vdd), .A(_16876_), .B(_16880_), .C(_16620_), .Y(_16887_) );
NAND3X1 NAND3X1_3826 ( .gnd(gnd), .vdd(vdd), .A(_16615_), .B(_16882_), .C(_16883_), .Y(_16888_) );
NAND3X1 NAND3X1_3827 ( .gnd(gnd), .vdd(vdd), .A(_16888_), .B(_16886_), .C(_16887_), .Y(_16889_) );
INVX1 INVX1_2372 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .Y(_16890_) );
OR2X2 OR2X2_396 ( .gnd(gnd), .vdd(vdd), .A(_16869_), .B(_16890_), .Y(_16891_) );
NAND2X1 NAND2X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_16890_), .B(_16869_), .Y(_16892_) );
NAND2X1 NAND2X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_16892_), .B(_16891_), .Y(_16893_) );
INVX2 INVX2_589 ( .gnd(gnd), .vdd(vdd), .A(_16893_), .Y(_16894_) );
XNOR2X1 XNOR2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_14972_), .B(_16894_), .Y(_16895_) );
NAND3X1 NAND3X1_3828 ( .gnd(gnd), .vdd(vdd), .A(_16895_), .B(_16889_), .C(_16885_), .Y(_16896_) );
AOI21X1 AOI21X1_2352 ( .gnd(gnd), .vdd(vdd), .A(_16888_), .B(_16887_), .C(_16886_), .Y(_13087_) );
AOI21X1 AOI21X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_16884_), .B(_16881_), .C(_16817_), .Y(_13088_) );
INVX1 INVX1_2373 ( .gnd(gnd), .vdd(vdd), .A(_16895_), .Y(_13089_) );
OAI21X1 OAI21X1_2687 ( .gnd(gnd), .vdd(vdd), .A(_13087_), .B(_13088_), .C(_13089_), .Y(_13090_) );
AOI21X1 AOI21X1_2354 ( .gnd(gnd), .vdd(vdd), .A(_16896_), .B(_13090_), .C(bloque_datos_36_bF_buf0_), .Y(_13091_) );
INVX1 INVX1_2374 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf3_), .Y(_13092_) );
NAND3X1 NAND3X1_3829 ( .gnd(gnd), .vdd(vdd), .A(_13089_), .B(_16889_), .C(_16885_), .Y(_13093_) );
OAI21X1 OAI21X1_2688 ( .gnd(gnd), .vdd(vdd), .A(_13087_), .B(_13088_), .C(_16895_), .Y(_13094_) );
AOI21X1 AOI21X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_13093_), .B(_13094_), .C(_13092_), .Y(_13095_) );
OAI21X1 OAI21X1_2689 ( .gnd(gnd), .vdd(vdd), .A(_13091_), .B(_13095_), .C(_16816_), .Y(_13096_) );
NAND3X1 NAND3X1_3830 ( .gnd(gnd), .vdd(vdd), .A(_13092_), .B(_13093_), .C(_13094_), .Y(_13097_) );
NAND3X1 NAND3X1_3831 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf2_), .B(_16896_), .C(_13090_), .Y(_13098_) );
NAND3X1 NAND3X1_3832 ( .gnd(gnd), .vdd(vdd), .A(_16634_), .B(_13097_), .C(_13098_), .Y(_13099_) );
NAND3X1 NAND3X1_3833 ( .gnd(gnd), .vdd(vdd), .A(_16815_), .B(_13099_), .C(_13096_), .Y(_13100_) );
OAI21X1 OAI21X1_2690 ( .gnd(gnd), .vdd(vdd), .A(_16579_), .B(_16637_), .C(_16633_), .Y(_13101_) );
OAI21X1 OAI21X1_2691 ( .gnd(gnd), .vdd(vdd), .A(_13091_), .B(_13095_), .C(_16634_), .Y(_13102_) );
NAND3X1 NAND3X1_3834 ( .gnd(gnd), .vdd(vdd), .A(_16816_), .B(_13097_), .C(_13098_), .Y(_13103_) );
NAND3X1 NAND3X1_3835 ( .gnd(gnd), .vdd(vdd), .A(_13101_), .B(_13103_), .C(_13102_), .Y(_13104_) );
NAND2X1 NAND2X1_2206 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf0_), .B(_16893_), .Y(_13105_) );
OR2X2 OR2X2_397 ( .gnd(gnd), .vdd(vdd), .A(_16893_), .B(bloque_datos_24_bF_buf4_), .Y(_13106_) );
NAND2X1 NAND2X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_13105_), .B(_13106_), .Y(_13107_) );
INVX2 INVX2_590 ( .gnd(gnd), .vdd(vdd), .A(_13107_), .Y(_13108_) );
XNOR2X1 XNOR2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_15002_), .B(_13108_), .Y(_13109_) );
NAND3X1 NAND3X1_3836 ( .gnd(gnd), .vdd(vdd), .A(_13109_), .B(_13100_), .C(_13104_), .Y(_13110_) );
AOI21X1 AOI21X1_2356 ( .gnd(gnd), .vdd(vdd), .A(_13103_), .B(_13102_), .C(_13101_), .Y(_13111_) );
AOI21X1 AOI21X1_2357 ( .gnd(gnd), .vdd(vdd), .A(_13099_), .B(_13096_), .C(_16815_), .Y(_13112_) );
INVX1 INVX1_2375 ( .gnd(gnd), .vdd(vdd), .A(_13109_), .Y(_13113_) );
OAI21X1 OAI21X1_2692 ( .gnd(gnd), .vdd(vdd), .A(_13111_), .B(_13112_), .C(_13113_), .Y(_13114_) );
AOI21X1 AOI21X1_2358 ( .gnd(gnd), .vdd(vdd), .A(_13110_), .B(_13114_), .C(bloque_datos_52_bF_buf1_), .Y(_13115_) );
INVX1 INVX1_2376 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf0_), .Y(_13116_) );
NAND3X1 NAND3X1_3837 ( .gnd(gnd), .vdd(vdd), .A(_13113_), .B(_13100_), .C(_13104_), .Y(_13117_) );
OAI21X1 OAI21X1_2693 ( .gnd(gnd), .vdd(vdd), .A(_13111_), .B(_13112_), .C(_13109_), .Y(_13118_) );
AOI21X1 AOI21X1_2359 ( .gnd(gnd), .vdd(vdd), .A(_13117_), .B(_13118_), .C(_13116_), .Y(_13119_) );
OAI21X1 OAI21X1_2694 ( .gnd(gnd), .vdd(vdd), .A(_13115_), .B(_13119_), .C(_16812_), .Y(_13120_) );
INVX2 INVX2_591 ( .gnd(gnd), .vdd(vdd), .A(_16812_), .Y(_13121_) );
NAND3X1 NAND3X1_3838 ( .gnd(gnd), .vdd(vdd), .A(_13116_), .B(_13117_), .C(_13118_), .Y(_13122_) );
NAND3X1 NAND3X1_3839 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf4_), .B(_13110_), .C(_13114_), .Y(_13123_) );
NAND3X1 NAND3X1_3840 ( .gnd(gnd), .vdd(vdd), .A(_13121_), .B(_13122_), .C(_13123_), .Y(_13124_) );
NAND3X1 NAND3X1_3841 ( .gnd(gnd), .vdd(vdd), .A(_13124_), .B(_16810_), .C(_13120_), .Y(_13125_) );
OAI21X1 OAI21X1_2695 ( .gnd(gnd), .vdd(vdd), .A(_16651_), .B(_16647_), .C(_16642_), .Y(_13126_) );
OAI21X1 OAI21X1_2696 ( .gnd(gnd), .vdd(vdd), .A(_13115_), .B(_13119_), .C(_13121_), .Y(_13127_) );
NAND3X1 NAND3X1_3842 ( .gnd(gnd), .vdd(vdd), .A(_16812_), .B(_13122_), .C(_13123_), .Y(_13128_) );
NAND3X1 NAND3X1_3843 ( .gnd(gnd), .vdd(vdd), .A(_13128_), .B(_13127_), .C(_13126_), .Y(_13129_) );
NAND2X1 NAND2X1_2208 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf0_), .B(_13107_), .Y(_13130_) );
OR2X2 OR2X2_398 ( .gnd(gnd), .vdd(vdd), .A(_13107_), .B(bloque_datos_40_bF_buf4_), .Y(_13131_) );
NAND2X1 NAND2X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_13130_), .B(_13131_), .Y(_13132_) );
INVX2 INVX2_592 ( .gnd(gnd), .vdd(vdd), .A(_13132_), .Y(_13133_) );
XNOR2X1 XNOR2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_13133_), .Y(_13134_) );
NAND3X1 NAND3X1_3844 ( .gnd(gnd), .vdd(vdd), .A(_13134_), .B(_13125_), .C(_13129_), .Y(_13135_) );
AOI21X1 AOI21X1_2360 ( .gnd(gnd), .vdd(vdd), .A(_13128_), .B(_13127_), .C(_13126_), .Y(_13136_) );
AOI21X1 AOI21X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_13124_), .B(_13120_), .C(_16810_), .Y(_13137_) );
INVX1 INVX1_2377 ( .gnd(gnd), .vdd(vdd), .A(_13134_), .Y(_13138_) );
OAI21X1 OAI21X1_2697 ( .gnd(gnd), .vdd(vdd), .A(_13136_), .B(_13137_), .C(_13138_), .Y(_13139_) );
AOI21X1 AOI21X1_2362 ( .gnd(gnd), .vdd(vdd), .A(_13135_), .B(_13139_), .C(bloque_datos_68_bF_buf0_), .Y(_13140_) );
INVX1 INVX1_2378 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf3_), .Y(_13141_) );
NAND3X1 NAND3X1_3845 ( .gnd(gnd), .vdd(vdd), .A(_13138_), .B(_13125_), .C(_13129_), .Y(_13142_) );
OAI21X1 OAI21X1_2698 ( .gnd(gnd), .vdd(vdd), .A(_13136_), .B(_13137_), .C(_13134_), .Y(_13143_) );
AOI21X1 AOI21X1_2363 ( .gnd(gnd), .vdd(vdd), .A(_13142_), .B(_13143_), .C(_13141_), .Y(_13144_) );
OAI21X1 OAI21X1_2699 ( .gnd(gnd), .vdd(vdd), .A(_13140_), .B(_13144_), .C(_16809_), .Y(_13145_) );
NAND3X1 NAND3X1_3846 ( .gnd(gnd), .vdd(vdd), .A(_13141_), .B(_13142_), .C(_13143_), .Y(_13146_) );
NAND3X1 NAND3X1_3847 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf2_), .B(_13135_), .C(_13139_), .Y(_13147_) );
NAND3X1 NAND3X1_3848 ( .gnd(gnd), .vdd(vdd), .A(_16658_), .B(_13146_), .C(_13147_), .Y(_13148_) );
NAND3X1 NAND3X1_3849 ( .gnd(gnd), .vdd(vdd), .A(_16808_), .B(_13148_), .C(_13145_), .Y(_13149_) );
INVX1 INVX1_2379 ( .gnd(gnd), .vdd(vdd), .A(_16576_), .Y(_13150_) );
AOI21X1 AOI21X1_2364 ( .gnd(gnd), .vdd(vdd), .A(_16653_), .B(_16656_), .C(_16445_), .Y(_13151_) );
OAI21X1 OAI21X1_2700 ( .gnd(gnd), .vdd(vdd), .A(_13151_), .B(_13150_), .C(_16657_), .Y(_13152_) );
OAI21X1 OAI21X1_2701 ( .gnd(gnd), .vdd(vdd), .A(_13140_), .B(_13144_), .C(_16658_), .Y(_13153_) );
NAND3X1 NAND3X1_3850 ( .gnd(gnd), .vdd(vdd), .A(_16809_), .B(_13146_), .C(_13147_), .Y(_13154_) );
NAND3X1 NAND3X1_3851 ( .gnd(gnd), .vdd(vdd), .A(_13152_), .B(_13154_), .C(_13153_), .Y(_13155_) );
NAND2X1 NAND2X1_2210 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf0_), .B(_13132_), .Y(_13156_) );
OR2X2 OR2X2_399 ( .gnd(gnd), .vdd(vdd), .A(_13132_), .B(bloque_datos_56_bF_buf4_), .Y(_13157_) );
NAND2X1 NAND2X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_13156_), .B(_13157_), .Y(_13158_) );
INVX2 INVX2_593 ( .gnd(gnd), .vdd(vdd), .A(_13158_), .Y(_13159_) );
XNOR2X1 XNOR2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_15068_), .B(_13159_), .Y(_13160_) );
NAND3X1 NAND3X1_3852 ( .gnd(gnd), .vdd(vdd), .A(_13160_), .B(_13149_), .C(_13155_), .Y(_13161_) );
AOI21X1 AOI21X1_2365 ( .gnd(gnd), .vdd(vdd), .A(_13154_), .B(_13153_), .C(_13152_), .Y(_13162_) );
AOI21X1 AOI21X1_2366 ( .gnd(gnd), .vdd(vdd), .A(_13148_), .B(_13145_), .C(_16808_), .Y(_13163_) );
INVX1 INVX1_2380 ( .gnd(gnd), .vdd(vdd), .A(_13160_), .Y(_13164_) );
OAI21X1 OAI21X1_2702 ( .gnd(gnd), .vdd(vdd), .A(_13162_), .B(_13163_), .C(_13164_), .Y(_13165_) );
AOI21X1 AOI21X1_2367 ( .gnd(gnd), .vdd(vdd), .A(_13161_), .B(_13165_), .C(bloque_datos_84_bF_buf1_), .Y(_13166_) );
INVX1 INVX1_2381 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf0_), .Y(_13167_) );
NAND3X1 NAND3X1_3853 ( .gnd(gnd), .vdd(vdd), .A(_13164_), .B(_13149_), .C(_13155_), .Y(_13168_) );
OAI21X1 OAI21X1_2703 ( .gnd(gnd), .vdd(vdd), .A(_13162_), .B(_13163_), .C(_13160_), .Y(_13169_) );
AOI21X1 AOI21X1_2368 ( .gnd(gnd), .vdd(vdd), .A(_13168_), .B(_13169_), .C(_13167_), .Y(_13170_) );
OAI21X1 OAI21X1_2704 ( .gnd(gnd), .vdd(vdd), .A(_13166_), .B(_13170_), .C(_16806_), .Y(_13171_) );
NAND3X1 NAND3X1_3854 ( .gnd(gnd), .vdd(vdd), .A(_13167_), .B(_13168_), .C(_13169_), .Y(_13172_) );
NAND3X1 NAND3X1_3855 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf4_), .B(_13161_), .C(_13165_), .Y(_13173_) );
NAND3X1 NAND3X1_3856 ( .gnd(gnd), .vdd(vdd), .A(_16670_), .B(_13172_), .C(_13173_), .Y(_13174_) );
NAND3X1 NAND3X1_3857 ( .gnd(gnd), .vdd(vdd), .A(_13171_), .B(_13174_), .C(_16805_), .Y(_13175_) );
NAND2X1 NAND2X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_16668_), .B(_16674_), .Y(_13176_) );
OAI21X1 OAI21X1_2705 ( .gnd(gnd), .vdd(vdd), .A(_13166_), .B(_13170_), .C(_16670_), .Y(_13177_) );
NAND3X1 NAND3X1_3858 ( .gnd(gnd), .vdd(vdd), .A(_16806_), .B(_13172_), .C(_13173_), .Y(_13178_) );
NAND3X1 NAND3X1_3859 ( .gnd(gnd), .vdd(vdd), .A(_13176_), .B(_13178_), .C(_13177_), .Y(_13179_) );
NOR2X1 NOR2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf1_), .B(_13159_), .Y(_13180_) );
NAND2X1 NAND2X1_2213 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf0_), .B(_13159_), .Y(_13181_) );
INVX1 INVX1_2382 ( .gnd(gnd), .vdd(vdd), .A(_13181_), .Y(_13182_) );
NOR2X1 NOR2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_13180_), .B(_13182_), .Y(_13183_) );
XOR2X1 XOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_15101_), .B(_13183_), .Y(_13184_) );
NAND3X1 NAND3X1_3860 ( .gnd(gnd), .vdd(vdd), .A(_13184_), .B(_13179_), .C(_13175_), .Y(_13185_) );
AOI21X1 AOI21X1_2369 ( .gnd(gnd), .vdd(vdd), .A(_13178_), .B(_13177_), .C(_13176_), .Y(_13186_) );
AOI21X1 AOI21X1_2370 ( .gnd(gnd), .vdd(vdd), .A(_13174_), .B(_13171_), .C(_16805_), .Y(_13187_) );
INVX1 INVX1_2383 ( .gnd(gnd), .vdd(vdd), .A(_13184_), .Y(_13188_) );
OAI21X1 OAI21X1_2706 ( .gnd(gnd), .vdd(vdd), .A(_13186_), .B(_13187_), .C(_13188_), .Y(_13189_) );
AOI21X1 AOI21X1_2371 ( .gnd(gnd), .vdd(vdd), .A(_13185_), .B(_13189_), .C(module_3_W_132_), .Y(_13190_) );
INVX1 INVX1_2384 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_132_), .Y(_13191_) );
NAND3X1 NAND3X1_3861 ( .gnd(gnd), .vdd(vdd), .A(_13188_), .B(_13179_), .C(_13175_), .Y(_13192_) );
OAI21X1 OAI21X1_2707 ( .gnd(gnd), .vdd(vdd), .A(_13186_), .B(_13187_), .C(_13184_), .Y(_13193_) );
AOI21X1 AOI21X1_2372 ( .gnd(gnd), .vdd(vdd), .A(_13192_), .B(_13193_), .C(_13191_), .Y(_13194_) );
OAI21X1 OAI21X1_2708 ( .gnd(gnd), .vdd(vdd), .A(_13190_), .B(_13194_), .C(_16676_), .Y(_13195_) );
INVX2 INVX2_594 ( .gnd(gnd), .vdd(vdd), .A(_16676_), .Y(_13196_) );
NAND3X1 NAND3X1_3862 ( .gnd(gnd), .vdd(vdd), .A(_13191_), .B(_13192_), .C(_13193_), .Y(_13197_) );
NAND3X1 NAND3X1_3863 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_132_), .B(_13185_), .C(_13189_), .Y(_13198_) );
NAND3X1 NAND3X1_3864 ( .gnd(gnd), .vdd(vdd), .A(_13196_), .B(_13197_), .C(_13198_), .Y(_13199_) );
AOI21X1 AOI21X1_2373 ( .gnd(gnd), .vdd(vdd), .A(_13199_), .B(_13195_), .C(_16804_), .Y(_13200_) );
AND2X2 AND2X2_379 ( .gnd(gnd), .vdd(vdd), .A(_16683_), .B(_16680_), .Y(_13201_) );
OAI21X1 OAI21X1_2709 ( .gnd(gnd), .vdd(vdd), .A(_13190_), .B(_13194_), .C(_13196_), .Y(_13202_) );
NAND3X1 NAND3X1_3865 ( .gnd(gnd), .vdd(vdd), .A(_16676_), .B(_13197_), .C(_13198_), .Y(_13203_) );
AOI21X1 AOI21X1_2374 ( .gnd(gnd), .vdd(vdd), .A(_13203_), .B(_13202_), .C(_13201_), .Y(_13204_) );
NAND2X1 NAND2X1_2214 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf2_), .B(_13183_), .Y(_13205_) );
OR2X2 OR2X2_400 ( .gnd(gnd), .vdd(vdd), .A(_13183_), .B(bloque_datos_88_bF_buf1_), .Y(_13206_) );
NAND2X1 NAND2X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_13205_), .B(_13206_), .Y(_13207_) );
OAI21X1 OAI21X1_2710 ( .gnd(gnd), .vdd(vdd), .A(_13200_), .B(_13204_), .C(_13207_), .Y(_13208_) );
AOI21X1 AOI21X1_2375 ( .gnd(gnd), .vdd(vdd), .A(_13197_), .B(_13198_), .C(_13196_), .Y(_13209_) );
NOR3X1 NOR3X1_503 ( .gnd(gnd), .vdd(vdd), .A(_13190_), .B(_16676_), .C(_13194_), .Y(_13210_) );
OAI21X1 OAI21X1_2711 ( .gnd(gnd), .vdd(vdd), .A(_13210_), .B(_13209_), .C(_13201_), .Y(_13211_) );
NAND3X1 NAND3X1_3866 ( .gnd(gnd), .vdd(vdd), .A(_16804_), .B(_13199_), .C(_13195_), .Y(_13212_) );
INVX2 INVX2_595 ( .gnd(gnd), .vdd(vdd), .A(_13207_), .Y(_13213_) );
NAND3X1 NAND3X1_3867 ( .gnd(gnd), .vdd(vdd), .A(_13212_), .B(_13213_), .C(_13211_), .Y(_13214_) );
NAND2X1 NAND2X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_13208_), .B(_13214_), .Y(_13215_) );
NAND3X1 NAND3X1_3868 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_148_), .B(_15134_), .C(_13215_), .Y(_13216_) );
INVX1 INVX1_2385 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_148_), .Y(_13217_) );
AOI21X1 AOI21X1_2376 ( .gnd(gnd), .vdd(vdd), .A(_13212_), .B(_13211_), .C(_13207_), .Y(_13218_) );
NAND2X1 NAND2X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_13212_), .B(_13211_), .Y(_13219_) );
OAI21X1 OAI21X1_2712 ( .gnd(gnd), .vdd(vdd), .A(_13219_), .B(_13213_), .C(_15134_), .Y(_13220_) );
OAI21X1 OAI21X1_2713 ( .gnd(gnd), .vdd(vdd), .A(_13220_), .B(_13218_), .C(_13217_), .Y(_13221_) );
AOI21X1 AOI21X1_2377 ( .gnd(gnd), .vdd(vdd), .A(_13216_), .B(_13221_), .C(_16689_), .Y(_13222_) );
OAI21X1 OAI21X1_2714 ( .gnd(gnd), .vdd(vdd), .A(_13220_), .B(_13218_), .C(module_3_W_148_), .Y(_13223_) );
NAND3X1 NAND3X1_3869 ( .gnd(gnd), .vdd(vdd), .A(_13217_), .B(_15134_), .C(_13215_), .Y(_13224_) );
AOI21X1 AOI21X1_2378 ( .gnd(gnd), .vdd(vdd), .A(_13224_), .B(_13223_), .C(_16688_), .Y(_13225_) );
OAI21X1 OAI21X1_2715 ( .gnd(gnd), .vdd(vdd), .A(_13225_), .B(_13222_), .C(_16803_), .Y(_13226_) );
NAND2X1 NAND2X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_16690_), .B(_16694_), .Y(_13227_) );
NAND3X1 NAND3X1_3870 ( .gnd(gnd), .vdd(vdd), .A(_16688_), .B(_13224_), .C(_13223_), .Y(_13228_) );
NAND3X1 NAND3X1_3871 ( .gnd(gnd), .vdd(vdd), .A(_16689_), .B(_13216_), .C(_13221_), .Y(_13229_) );
NAND3X1 NAND3X1_3872 ( .gnd(gnd), .vdd(vdd), .A(_13227_), .B(_13228_), .C(_13229_), .Y(_13230_) );
NAND2X1 NAND2X1_2219 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_136_), .B(_13207_), .Y(_13231_) );
OR2X2 OR2X2_401 ( .gnd(gnd), .vdd(vdd), .A(_13207_), .B(module_3_W_136_), .Y(_13232_) );
NAND2X1 NAND2X1_2220 ( .gnd(gnd), .vdd(vdd), .A(_13231_), .B(_13232_), .Y(_13233_) );
NAND3X1 NAND3X1_3873 ( .gnd(gnd), .vdd(vdd), .A(_13230_), .B(_13233_), .C(_13226_), .Y(_13234_) );
NAND2X1 NAND2X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_13230_), .B(_13226_), .Y(_13235_) );
INVX2 INVX2_596 ( .gnd(gnd), .vdd(vdd), .A(_13233_), .Y(_13236_) );
AOI21X1 AOI21X1_2379 ( .gnd(gnd), .vdd(vdd), .A(_13236_), .B(_13235_), .C(_15419_), .Y(_13237_) );
NAND3X1 NAND3X1_3874 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_164_), .B(_13234_), .C(_13237_), .Y(_13238_) );
INVX1 INVX1_2386 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_164_), .Y(_13239_) );
AOI21X1 AOI21X1_2380 ( .gnd(gnd), .vdd(vdd), .A(_13228_), .B(_13229_), .C(_13227_), .Y(_13240_) );
NAND3X1 NAND3X1_3875 ( .gnd(gnd), .vdd(vdd), .A(_16688_), .B(_13216_), .C(_13221_), .Y(_13241_) );
NAND3X1 NAND3X1_3876 ( .gnd(gnd), .vdd(vdd), .A(_16689_), .B(_13224_), .C(_13223_), .Y(_13242_) );
AOI21X1 AOI21X1_2381 ( .gnd(gnd), .vdd(vdd), .A(_13241_), .B(_13242_), .C(_16803_), .Y(_13243_) );
OAI21X1 OAI21X1_2716 ( .gnd(gnd), .vdd(vdd), .A(_13240_), .B(_13243_), .C(_13236_), .Y(_13244_) );
NAND3X1 NAND3X1_3877 ( .gnd(gnd), .vdd(vdd), .A(_15167_), .B(_13234_), .C(_13244_), .Y(_13245_) );
NAND2X1 NAND2X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_13239_), .B(_13245_), .Y(_13246_) );
AOI21X1 AOI21X1_2382 ( .gnd(gnd), .vdd(vdd), .A(_13246_), .B(_13238_), .C(_16699_), .Y(_13247_) );
INVX1 INVX1_2387 ( .gnd(gnd), .vdd(vdd), .A(_16699_), .Y(_13248_) );
NAND2X1 NAND2X1_2223 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_164_), .B(_13245_), .Y(_13249_) );
NAND3X1 NAND3X1_3878 ( .gnd(gnd), .vdd(vdd), .A(_13239_), .B(_13234_), .C(_13237_), .Y(_13250_) );
AOI21X1 AOI21X1_2383 ( .gnd(gnd), .vdd(vdd), .A(_13249_), .B(_13250_), .C(_13248_), .Y(_13251_) );
OAI21X1 OAI21X1_2717 ( .gnd(gnd), .vdd(vdd), .A(_13251_), .B(_13247_), .C(_16802_), .Y(_13252_) );
NAND3X1 NAND3X1_3879 ( .gnd(gnd), .vdd(vdd), .A(_13248_), .B(_13249_), .C(_13250_), .Y(_13253_) );
NAND3X1 NAND3X1_3880 ( .gnd(gnd), .vdd(vdd), .A(_16699_), .B(_13246_), .C(_13238_), .Y(_13254_) );
NAND3X1 NAND3X1_3881 ( .gnd(gnd), .vdd(vdd), .A(_16801_), .B(_13253_), .C(_13254_), .Y(_13255_) );
NAND2X1 NAND2X1_2224 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_152_), .B(_13233_), .Y(_13256_) );
OR2X2 OR2X2_402 ( .gnd(gnd), .vdd(vdd), .A(_13233_), .B(module_3_W_152_), .Y(_13257_) );
NAND2X1 NAND2X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_13256_), .B(_13257_), .Y(_13258_) );
NAND3X1 NAND3X1_3882 ( .gnd(gnd), .vdd(vdd), .A(_13255_), .B(_13258_), .C(_13252_), .Y(_13259_) );
AOI21X1 AOI21X1_2384 ( .gnd(gnd), .vdd(vdd), .A(_13255_), .B(_13252_), .C(_13258_), .Y(_13260_) );
NOR2X1 NOR2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_15397_), .B(_13260_), .Y(_13261_) );
NAND3X1 NAND3X1_3883 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_180_), .B(_13259_), .C(_13261_), .Y(_13262_) );
INVX1 INVX1_2388 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_180_), .Y(_13263_) );
NAND2X1 NAND2X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_15200_), .B(_13259_), .Y(_13264_) );
OAI21X1 OAI21X1_2718 ( .gnd(gnd), .vdd(vdd), .A(_13264_), .B(_13260_), .C(_13263_), .Y(_13265_) );
AOI21X1 AOI21X1_2385 ( .gnd(gnd), .vdd(vdd), .A(_13265_), .B(_13262_), .C(_16712_), .Y(_13266_) );
OAI21X1 OAI21X1_2719 ( .gnd(gnd), .vdd(vdd), .A(_13264_), .B(_13260_), .C(module_3_W_180_), .Y(_13267_) );
NAND3X1 NAND3X1_3884 ( .gnd(gnd), .vdd(vdd), .A(_13263_), .B(_13259_), .C(_13261_), .Y(_13268_) );
AOI21X1 AOI21X1_2386 ( .gnd(gnd), .vdd(vdd), .A(_13267_), .B(_13268_), .C(_16711_), .Y(_13269_) );
OAI21X1 OAI21X1_2720 ( .gnd(gnd), .vdd(vdd), .A(_13269_), .B(_13266_), .C(_16799_), .Y(_13270_) );
OAI21X1 OAI21X1_2721 ( .gnd(gnd), .vdd(vdd), .A(_16719_), .B(_16566_), .C(_16713_), .Y(_13271_) );
NAND3X1 NAND3X1_3885 ( .gnd(gnd), .vdd(vdd), .A(_16711_), .B(_13267_), .C(_13268_), .Y(_13272_) );
NAND3X1 NAND3X1_3886 ( .gnd(gnd), .vdd(vdd), .A(_16712_), .B(_13265_), .C(_13262_), .Y(_13273_) );
NAND3X1 NAND3X1_3887 ( .gnd(gnd), .vdd(vdd), .A(_13272_), .B(_13271_), .C(_13273_), .Y(_13274_) );
NAND2X1 NAND2X1_2227 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_168_), .B(_13258_), .Y(_13275_) );
OR2X2 OR2X2_403 ( .gnd(gnd), .vdd(vdd), .A(_13258_), .B(module_3_W_168_), .Y(_13276_) );
NAND2X1 NAND2X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_13275_), .B(_13276_), .Y(_13277_) );
NAND3X1 NAND3X1_3888 ( .gnd(gnd), .vdd(vdd), .A(_13274_), .B(_13277_), .C(_13270_), .Y(_13278_) );
NAND2X1 NAND2X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_13274_), .B(_13270_), .Y(_13279_) );
INVX2 INVX2_597 ( .gnd(gnd), .vdd(vdd), .A(_13277_), .Y(_13280_) );
AOI21X1 AOI21X1_2387 ( .gnd(gnd), .vdd(vdd), .A(_13280_), .B(_13279_), .C(_15364_), .Y(_13281_) );
NAND3X1 NAND3X1_3889 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_196_), .B(_13278_), .C(_13281_), .Y(_13282_) );
INVX1 INVX1_2389 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_196_), .Y(_13283_) );
AOI21X1 AOI21X1_2388 ( .gnd(gnd), .vdd(vdd), .A(_13272_), .B(_13273_), .C(_13271_), .Y(_13284_) );
NOR3X1 NOR3X1_504 ( .gnd(gnd), .vdd(vdd), .A(_13266_), .B(_16799_), .C(_13269_), .Y(_13285_) );
OAI21X1 OAI21X1_2722 ( .gnd(gnd), .vdd(vdd), .A(_13285_), .B(_13284_), .C(_13280_), .Y(_13286_) );
NAND3X1 NAND3X1_3890 ( .gnd(gnd), .vdd(vdd), .A(_15233_), .B(_13278_), .C(_13286_), .Y(_13287_) );
NAND2X1 NAND2X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_13283_), .B(_13287_), .Y(_13288_) );
AOI21X1 AOI21X1_2389 ( .gnd(gnd), .vdd(vdd), .A(_13282_), .B(_13288_), .C(_16724_), .Y(_13289_) );
INVX1 INVX1_2390 ( .gnd(gnd), .vdd(vdd), .A(_16717_), .Y(_13290_) );
NAND2X1 NAND2X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_16720_), .B(_13290_), .Y(_13291_) );
NOR2X1 NOR2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_16565_), .B(_13291_), .Y(_13292_) );
NAND2X1 NAND2X1_2232 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_196_), .B(_13287_), .Y(_13293_) );
NAND3X1 NAND3X1_3891 ( .gnd(gnd), .vdd(vdd), .A(_13283_), .B(_13278_), .C(_13281_), .Y(_13294_) );
AOI21X1 AOI21X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_13294_), .B(_13293_), .C(_13292_), .Y(_13295_) );
OAI21X1 OAI21X1_2723 ( .gnd(gnd), .vdd(vdd), .A(_13289_), .B(_13295_), .C(_16797_), .Y(_13296_) );
OAI21X1 OAI21X1_2724 ( .gnd(gnd), .vdd(vdd), .A(_16727_), .B(_16563_), .C(_16726_), .Y(_13297_) );
NAND3X1 NAND3X1_3892 ( .gnd(gnd), .vdd(vdd), .A(_13292_), .B(_13294_), .C(_13293_), .Y(_13298_) );
NAND3X1 NAND3X1_3893 ( .gnd(gnd), .vdd(vdd), .A(_16724_), .B(_13282_), .C(_13288_), .Y(_13299_) );
NAND3X1 NAND3X1_3894 ( .gnd(gnd), .vdd(vdd), .A(_13298_), .B(_13299_), .C(_13297_), .Y(_13300_) );
NAND2X1 NAND2X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_13300_), .B(_13296_), .Y(_13301_) );
NAND2X1 NAND2X1_2234 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_184_), .B(_13277_), .Y(_13302_) );
OR2X2 OR2X2_404 ( .gnd(gnd), .vdd(vdd), .A(_13277_), .B(module_3_W_184_), .Y(_13303_) );
NAND2X1 NAND2X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_13302_), .B(_13303_), .Y(_13304_) );
INVX2 INVX2_598 ( .gnd(gnd), .vdd(vdd), .A(_13304_), .Y(_13305_) );
OR2X2 OR2X2_405 ( .gnd(gnd), .vdd(vdd), .A(_13301_), .B(_13305_), .Y(_13306_) );
AOI21X1 AOI21X1_2391 ( .gnd(gnd), .vdd(vdd), .A(_13300_), .B(_13296_), .C(_13304_), .Y(_13307_) );
NOR2X1 NOR2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_15343_), .B(_13307_), .Y(_13308_) );
NAND3X1 NAND3X1_3895 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_212_), .B(_13306_), .C(_13308_), .Y(_13309_) );
INVX1 INVX1_2391 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_212_), .Y(_13310_) );
OAI21X1 OAI21X1_2725 ( .gnd(gnd), .vdd(vdd), .A(_13301_), .B(_13305_), .C(_15266_), .Y(_13311_) );
OAI21X1 OAI21X1_2726 ( .gnd(gnd), .vdd(vdd), .A(_13311_), .B(_13307_), .C(_13310_), .Y(_13312_) );
AOI21X1 AOI21X1_2392 ( .gnd(gnd), .vdd(vdd), .A(_13312_), .B(_13309_), .C(_16742_), .Y(_13313_) );
OAI21X1 OAI21X1_2727 ( .gnd(gnd), .vdd(vdd), .A(_13311_), .B(_13307_), .C(module_3_W_212_), .Y(_13314_) );
NAND3X1 NAND3X1_3896 ( .gnd(gnd), .vdd(vdd), .A(_13310_), .B(_13306_), .C(_13308_), .Y(_13315_) );
AOI21X1 AOI21X1_2393 ( .gnd(gnd), .vdd(vdd), .A(_13314_), .B(_13315_), .C(_16739_), .Y(_13316_) );
OAI21X1 OAI21X1_2728 ( .gnd(gnd), .vdd(vdd), .A(_13313_), .B(_13316_), .C(_16795_), .Y(_13317_) );
NAND3X1 NAND3X1_3897 ( .gnd(gnd), .vdd(vdd), .A(_16520_), .B(_16734_), .C(_16742_), .Y(_13318_) );
OAI21X1 OAI21X1_2729 ( .gnd(gnd), .vdd(vdd), .A(_16746_), .B(_16743_), .C(_13318_), .Y(_13319_) );
NAND3X1 NAND3X1_3898 ( .gnd(gnd), .vdd(vdd), .A(_16739_), .B(_13314_), .C(_13315_), .Y(_13320_) );
NAND3X1 NAND3X1_3899 ( .gnd(gnd), .vdd(vdd), .A(_16742_), .B(_13312_), .C(_13309_), .Y(_13321_) );
INVX1 INVX1_2392 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_0_), .Y(_17077_) );
INVX4 INVX4_15 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .Y(_17078_) );
NAND2X1 NAND2X1_2236 ( .gnd(gnd), .vdd(vdd), .A(nonce_iniciales[96]), .B(_17078_), .Y(_16898_) );
OAI21X1 OAI21X1_2730 ( .gnd(gnd), .vdd(vdd), .A(_17077_), .B(_17078_), .C(_16898_), .Y(_16897__0_) );
INVX1 INVX1_2393 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_1_), .Y(_16899_) );
NAND2X1 NAND2X1_2237 ( .gnd(gnd), .vdd(vdd), .A(nonce_iniciales[97]), .B(_17078_), .Y(_16900_) );
OAI21X1 OAI21X1_2731 ( .gnd(gnd), .vdd(vdd), .A(_17078_), .B(_16899_), .C(_16900_), .Y(_16897__1_) );
NAND2X1 NAND2X1_2238 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_5_), .B(module_3_W_4_), .Y(_16901_) );
NAND2X1 NAND2X1_2239 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_7_), .B(module_3_W_6_), .Y(_16902_) );
NOR2X1 NOR2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_16901_), .B(_16902_), .Y(_16903_) );
NAND2X1 NAND2X1_2240 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_25_), .B(module_3_W_24_), .Y(_16904_) );
NAND2X1 NAND2X1_2241 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_27_), .B(module_3_W_26_), .Y(_16905_) );
NOR2X1 NOR2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_16904_), .B(_16905_), .Y(_16906_) );
INVX1 INVX1_2394 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_2_), .Y(_16907_) );
OAI21X1 OAI21X1_2732 ( .gnd(gnd), .vdd(vdd), .A(_17077_), .B(_16899_), .C(_16907_), .Y(_16908_) );
NAND3X1 NAND3X1_3900 ( .gnd(gnd), .vdd(vdd), .A(_16908_), .B(_16903_), .C(_16906_), .Y(_16909_) );
INVX1 INVX1_2395 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_29_), .Y(_16910_) );
INVX1 INVX1_2396 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_28_), .Y(_16911_) );
NOR2X1 NOR2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_16910_), .B(_16911_), .Y(_16912_) );
INVX1 INVX1_2397 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_31_), .Y(_16913_) );
INVX1 INVX1_2398 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_30_), .Y(_16914_) );
NOR2X1 NOR2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_16913_), .B(_16914_), .Y(_16915_) );
NAND3X1 NAND3X1_3901 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_3_), .B(_16912_), .C(_16915_), .Y(_16916_) );
NOR2X1 NOR2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_16916_), .B(_16909_), .Y(_16917_) );
NAND2X1 NAND2X1_2242 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_17_), .B(module_3_W_16_), .Y(_16918_) );
NAND2X1 NAND2X1_2243 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_19_), .B(module_3_W_18_), .Y(_16919_) );
NOR2X1 NOR2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_16918_), .B(_16919_), .Y(_16920_) );
NAND2X1 NAND2X1_2244 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_22_), .B(module_3_W_21_), .Y(_16921_) );
NAND2X1 NAND2X1_2245 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_23_), .B(module_3_W_20_), .Y(_16922_) );
NOR2X1 NOR2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_16921_), .B(_16922_), .Y(_16923_) );
NAND2X1 NAND2X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_16920_), .B(_16923_), .Y(_16924_) );
NAND2X1 NAND2X1_2247 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_9_), .B(module_3_W_8_), .Y(_16925_) );
NAND2X1 NAND2X1_2248 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_11_), .B(module_3_W_10_), .Y(_16926_) );
NOR2X1 NOR2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_16925_), .B(_16926_), .Y(_16927_) );
NAND2X1 NAND2X1_2249 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_15_), .B(module_3_W_14_), .Y(_16928_) );
NAND2X1 NAND2X1_2250 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_13_), .B(module_3_W_12_), .Y(_16929_) );
NOR2X1 NOR2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_16928_), .B(_16929_), .Y(_16930_) );
NAND2X1 NAND2X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_16927_), .B(_16930_), .Y(_16931_) );
NOR2X1 NOR2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_16924_), .B(_16931_), .Y(_16932_) );
AOI21X1 AOI21X1_2394 ( .gnd(gnd), .vdd(vdd), .A(_16932_), .B(_16917_), .C(_17078_), .Y(_16933_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_2_), .B(nonce_iniciales[98]), .S(inicio_bF_buf6), .Y(_16934_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_2_), .B(_16934_), .S(_16933__bF_buf3), .Y(_16897__2_) );
NAND2X1 NAND2X1_2252 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_2_), .B(module_3_W_3_), .Y(_16935_) );
INVX1 INVX1_2399 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_3_), .Y(_16936_) );
NAND2X1 NAND2X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_16907_), .B(_16936_), .Y(_16937_) );
NAND2X1 NAND2X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_16935_), .B(_16937_), .Y(_16938_) );
NOR2X1 NOR2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf6), .B(nonce_iniciales[99]), .Y(_16939_) );
AOI21X1 AOI21X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_16938_), .B(_16933__bF_buf3), .C(_16939_), .Y(_16897__3_) );
XOR2X1 XOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_16935_), .B(module_3_W_4_), .Y(_16940_) );
NOR2X1 NOR2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[100]), .Y(_16941_) );
AOI21X1 AOI21X1_2396 ( .gnd(gnd), .vdd(vdd), .A(_16940_), .B(_16933__bF_buf3), .C(_16941_), .Y(_16897__4_) );
AND2X2 AND2X2_380 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_2_), .B(module_3_W_3_), .Y(_16942_) );
NAND2X1 NAND2X1_2255 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_4_), .B(_16942_), .Y(_16943_) );
XOR2X1 XOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_16943_), .B(module_3_W_5_), .Y(_16944_) );
NOR2X1 NOR2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf6), .B(nonce_iniciales[101]), .Y(_16945_) );
AOI21X1 AOI21X1_2397 ( .gnd(gnd), .vdd(vdd), .A(_16944_), .B(_16933__bF_buf0), .C(_16945_), .Y(_16897__5_) );
NOR2X1 NOR2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_16901_), .B(_16935_), .Y(_16946_) );
XNOR2X1 XNOR2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_16946_), .B(module_3_W_6_), .Y(_16947_) );
NOR2X1 NOR2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf6), .B(nonce_iniciales[102]), .Y(_16948_) );
AOI21X1 AOI21X1_2398 ( .gnd(gnd), .vdd(vdd), .A(_16947_), .B(_16933__bF_buf3), .C(_16948_), .Y(_16897__6_) );
NOR2X1 NOR2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[103]), .Y(_16949_) );
NAND2X1 NAND2X1_2256 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_6_), .B(_16946_), .Y(_16950_) );
XOR2X1 XOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_16950_), .B(module_3_W_7_), .Y(_16951_) );
AOI21X1 AOI21X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_16951_), .B(_16933__bF_buf3), .C(_16949_), .Y(_16897__7_) );
NOR3X1 NOR3X1_505 ( .gnd(gnd), .vdd(vdd), .A(_16901_), .B(_16902_), .C(_16935_), .Y(_16952_) );
XNOR2X1 XNOR2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_16952_), .B(module_3_W_8_), .Y(_16953_) );
NOR2X1 NOR2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[104]), .Y(_16954_) );
AOI21X1 AOI21X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_16953_), .B(_16933__bF_buf0), .C(_16954_), .Y(_16897__8_) );
AND2X2 AND2X2_381 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_5_), .B(module_3_W_4_), .Y(_16955_) );
AND2X2 AND2X2_382 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_7_), .B(module_3_W_6_), .Y(_16956_) );
NAND3X1 NAND3X1_3902 ( .gnd(gnd), .vdd(vdd), .A(_16955_), .B(_16956_), .C(_16942_), .Y(_16957_) );
INVX1 INVX1_2400 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_9_), .Y(_16958_) );
INVX1 INVX1_2401 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_8_), .Y(_16959_) );
OAI21X1 OAI21X1_2733 ( .gnd(gnd), .vdd(vdd), .A(_16957_), .B(_16959_), .C(_16958_), .Y(_16960_) );
OAI21X1 OAI21X1_2734 ( .gnd(gnd), .vdd(vdd), .A(_16925_), .B(_16957_), .C(_16960_), .Y(_16961_) );
NOR2X1 NOR2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[105]), .Y(_16962_) );
AOI21X1 AOI21X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_16961_), .B(_16933__bF_buf3), .C(_16962_), .Y(_16897__9_) );
NOR2X1 NOR2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_16925_), .B(_16957_), .Y(_16963_) );
XNOR2X1 XNOR2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_16963_), .B(module_3_W_10_), .Y(_16964_) );
NOR2X1 NOR2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[106]), .Y(_16965_) );
AOI21X1 AOI21X1_2402 ( .gnd(gnd), .vdd(vdd), .A(_16964_), .B(_16933__bF_buf1), .C(_16965_), .Y(_16897__10_) );
NOR2X1 NOR2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[107]), .Y(_16966_) );
NAND2X1 NAND2X1_2257 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_10_), .B(_16963_), .Y(_16967_) );
OR2X2 OR2X2_406 ( .gnd(gnd), .vdd(vdd), .A(_16967_), .B(module_3_W_11_), .Y(_16968_) );
NAND2X1 NAND2X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_16932_), .B(_16917_), .Y(_16969_) );
NAND2X1 NAND2X1_2259 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .B(_16969_), .Y(_16970_) );
AOI21X1 AOI21X1_2403 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_11_), .B(_16967_), .C(_16970_), .Y(_16971_) );
AOI21X1 AOI21X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_16968_), .B(_16971_), .C(_16966_), .Y(_16897__11_) );
INVX2 INVX2_599 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_12_), .Y(_16972_) );
NAND2X1 NAND2X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_16927_), .B(_16952_), .Y(_16973_) );
XNOR2X1 XNOR2X1_442 ( .gnd(gnd), .vdd(vdd), .A(_16973_), .B(_16972_), .Y(_16974_) );
NOR2X1 NOR2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .B(nonce_iniciales[108]), .Y(_16975_) );
AOI21X1 AOI21X1_2405 ( .gnd(gnd), .vdd(vdd), .A(_16974_), .B(_16933__bF_buf1), .C(_16975_), .Y(_16897__12_) );
NOR2X1 NOR2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf1), .B(nonce_iniciales[109]), .Y(_16976_) );
INVX1 INVX1_2402 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_13_), .Y(_16977_) );
NAND3X1 NAND3X1_3903 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_11_), .B(module_3_W_10_), .C(_16963_), .Y(_16978_) );
NOR2X1 NOR2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_16972_), .B(_16978_), .Y(_16979_) );
NAND2X1 NAND2X1_2261 ( .gnd(gnd), .vdd(vdd), .A(_16977_), .B(_16979_), .Y(_16980_) );
OAI21X1 OAI21X1_2735 ( .gnd(gnd), .vdd(vdd), .A(_16973_), .B(_16972_), .C(module_3_W_13_), .Y(_16981_) );
AND2X2 AND2X2_383 ( .gnd(gnd), .vdd(vdd), .A(_16933__bF_buf2), .B(_16981_), .Y(_16982_) );
AOI21X1 AOI21X1_2406 ( .gnd(gnd), .vdd(vdd), .A(_16980_), .B(_16982_), .C(_16976_), .Y(_16897__13_) );
INVX2 INVX2_600 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_14_), .Y(_16983_) );
OR2X2 OR2X2_407 ( .gnd(gnd), .vdd(vdd), .A(_16973_), .B(_16929_), .Y(_16984_) );
XNOR2X1 XNOR2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_16984_), .B(_16983_), .Y(_16985_) );
NOR2X1 NOR2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .B(nonce_iniciales[110]), .Y(_16986_) );
AOI21X1 AOI21X1_2407 ( .gnd(gnd), .vdd(vdd), .A(_16933__bF_buf1), .B(_16985_), .C(_16986_), .Y(_16897__14_) );
NOR2X1 NOR2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .B(nonce_iniciales[111]), .Y(_16987_) );
INVX1 INVX1_2403 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_15_), .Y(_16988_) );
NOR2X1 NOR2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_16929_), .B(_16978_), .Y(_16989_) );
NAND3X1 NAND3X1_3904 ( .gnd(gnd), .vdd(vdd), .A(_16988_), .B(module_3_W_14_), .C(_16989_), .Y(_16990_) );
OAI21X1 OAI21X1_2736 ( .gnd(gnd), .vdd(vdd), .A(_16984_), .B(_16983_), .C(module_3_W_15_), .Y(_16991_) );
AND2X2 AND2X2_384 ( .gnd(gnd), .vdd(vdd), .A(_16991_), .B(_16933__bF_buf1), .Y(_16992_) );
AOI21X1 AOI21X1_2408 ( .gnd(gnd), .vdd(vdd), .A(_16990_), .B(_16992_), .C(_16987_), .Y(_16897__15_) );
OR2X2 OR2X2_408 ( .gnd(gnd), .vdd(vdd), .A(_16925_), .B(_16926_), .Y(_16993_) );
OR2X2 OR2X2_409 ( .gnd(gnd), .vdd(vdd), .A(_16928_), .B(_16929_), .Y(_16994_) );
NOR3X1 NOR3X1_506 ( .gnd(gnd), .vdd(vdd), .A(_16994_), .B(_16993_), .C(_16957_), .Y(_16995_) );
NAND2X1 NAND2X1_2262 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_16_), .B(_16995_), .Y(_16996_) );
INVX1 INVX1_2404 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_16_), .Y(_16997_) );
OAI21X1 OAI21X1_2737 ( .gnd(gnd), .vdd(vdd), .A(_16931_), .B(_16957_), .C(_16997_), .Y(_16998_) );
NAND2X1 NAND2X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_16998_), .B(_16996_), .Y(_16999_) );
NOR2X1 NOR2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[112]), .Y(_17000_) );
AOI21X1 AOI21X1_2409 ( .gnd(gnd), .vdd(vdd), .A(_16933__bF_buf0), .B(_16999_), .C(_17000_), .Y(_16897__16_) );
NAND3X1 NAND3X1_3905 ( .gnd(gnd), .vdd(vdd), .A(_16927_), .B(_16930_), .C(_16952_), .Y(_17001_) );
NOR2X1 NOR2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_16997_), .B(_17001_), .Y(_17002_) );
XNOR2X1 XNOR2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_17002_), .B(module_3_W_17_), .Y(_17003_) );
NOR2X1 NOR2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[113]), .Y(_17004_) );
AOI21X1 AOI21X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_16933__bF_buf1), .B(_17003_), .C(_17004_), .Y(_16897__17_) );
INVX1 INVX1_2405 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_18_), .Y(_17005_) );
INVX1 INVX1_2406 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_17_), .Y(_17006_) );
OAI21X1 OAI21X1_2738 ( .gnd(gnd), .vdd(vdd), .A(_16996_), .B(_17006_), .C(_17005_), .Y(_17007_) );
NAND3X1 NAND3X1_3906 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_18_), .B(module_3_W_17_), .C(_17002_), .Y(_17008_) );
NAND2X1 NAND2X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_17008_), .B(_17007_), .Y(_17009_) );
NOR2X1 NOR2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .B(nonce_iniciales[114]), .Y(_17010_) );
AOI21X1 AOI21X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_16933__bF_buf2), .B(_17009_), .C(_17010_), .Y(_16897__18_) );
NOR2X1 NOR2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[115]), .Y(_17011_) );
OR2X2 OR2X2_410 ( .gnd(gnd), .vdd(vdd), .A(_17008_), .B(module_3_W_19_), .Y(_17012_) );
AOI21X1 AOI21X1_2412 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_19_), .B(_17008_), .C(_16970_), .Y(_17013_) );
AOI21X1 AOI21X1_2413 ( .gnd(gnd), .vdd(vdd), .A(_17012_), .B(_17013_), .C(_17011_), .Y(_16897__19_) );
INVX1 INVX1_2407 ( .gnd(gnd), .vdd(vdd), .A(_16920_), .Y(_17014_) );
NOR2X1 NOR2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_17014_), .B(_17001_), .Y(_17015_) );
NAND2X1 NAND2X1_2265 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_20_), .B(_17015_), .Y(_17016_) );
INVX2 INVX2_601 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_20_), .Y(_17017_) );
OAI21X1 OAI21X1_2739 ( .gnd(gnd), .vdd(vdd), .A(_17001_), .B(_17014_), .C(_17017_), .Y(_17018_) );
NAND2X1 NAND2X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_17018_), .B(_17016_), .Y(_17019_) );
NOR2X1 NOR2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .B(nonce_iniciales[116]), .Y(_17020_) );
AOI21X1 AOI21X1_2414 ( .gnd(gnd), .vdd(vdd), .A(_16933__bF_buf2), .B(_17019_), .C(_17020_), .Y(_16897__20_) );
INVX1 INVX1_2408 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_21_), .Y(_17021_) );
INVX1 INVX1_2409 ( .gnd(gnd), .vdd(vdd), .A(_16969_), .Y(_17022_) );
NAND2X1 NAND2X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_16920_), .B(_16995_), .Y(_17023_) );
NOR2X1 NOR2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_17017_), .B(_17023_), .Y(_17024_) );
AOI21X1 AOI21X1_2415 ( .gnd(gnd), .vdd(vdd), .A(_17021_), .B(_17024_), .C(_17022_), .Y(_17025_) );
AOI21X1 AOI21X1_2416 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_21_), .B(_17016_), .C(_17078_), .Y(_17026_) );
NOR2X1 NOR2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .B(nonce_iniciales[117]), .Y(_17027_) );
AOI21X1 AOI21X1_2417 ( .gnd(gnd), .vdd(vdd), .A(_17026_), .B(_17025_), .C(_17027_), .Y(_16897__21_) );
NOR2X1 NOR2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_17021_), .B(_17017_), .Y(_17028_) );
INVX1 INVX1_2410 ( .gnd(gnd), .vdd(vdd), .A(_17028_), .Y(_17029_) );
OAI21X1 OAI21X1_2740 ( .gnd(gnd), .vdd(vdd), .A(_17023_), .B(_17029_), .C(module_3_W_22_), .Y(_17030_) );
INVX1 INVX1_2411 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_22_), .Y(_17031_) );
NAND3X1 NAND3X1_3907 ( .gnd(gnd), .vdd(vdd), .A(_17031_), .B(_17028_), .C(_17015_), .Y(_17032_) );
AND2X2 AND2X2_385 ( .gnd(gnd), .vdd(vdd), .A(_17030_), .B(_17032_), .Y(_17033_) );
NOR2X1 NOR2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf1), .B(nonce_iniciales[118]), .Y(_17034_) );
AOI21X1 AOI21X1_2418 ( .gnd(gnd), .vdd(vdd), .A(_16933__bF_buf2), .B(_17033_), .C(_17034_), .Y(_16897__22_) );
NOR2X1 NOR2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .B(nonce_iniciales[119]), .Y(_17035_) );
INVX1 INVX1_2412 ( .gnd(gnd), .vdd(vdd), .A(_16921_), .Y(_17036_) );
NAND3X1 NAND3X1_3908 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_20_), .B(_17036_), .C(_17015_), .Y(_17037_) );
OR2X2 OR2X2_411 ( .gnd(gnd), .vdd(vdd), .A(_17037_), .B(module_3_W_23_), .Y(_17038_) );
AOI21X1 AOI21X1_2419 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_23_), .B(_17037_), .C(_16970_), .Y(_17039_) );
AOI21X1 AOI21X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_17038_), .B(_17039_), .C(_17035_), .Y(_16897__23_) );
NOR2X1 NOR2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_16924_), .B(_17001_), .Y(_17040_) );
XNOR2X1 XNOR2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_17040_), .B(module_3_W_24_), .Y(_17041_) );
NOR2X1 NOR2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .B(nonce_iniciales[120]), .Y(_17042_) );
AOI21X1 AOI21X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_16933__bF_buf2), .B(_17041_), .C(_17042_), .Y(_16897__24_) );
INVX1 INVX1_2413 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_25_), .Y(_17043_) );
AND2X2 AND2X2_386 ( .gnd(gnd), .vdd(vdd), .A(_17040_), .B(module_3_W_24_), .Y(_17044_) );
AOI21X1 AOI21X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_17043_), .B(_17044_), .C(_17022_), .Y(_17045_) );
NAND2X1 NAND2X1_2268 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_24_), .B(_17040_), .Y(_17046_) );
AOI21X1 AOI21X1_2423 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_25_), .B(_17046_), .C(_17078_), .Y(_17047_) );
NOR2X1 NOR2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .B(nonce_iniciales[121]), .Y(_17048_) );
AOI21X1 AOI21X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_17047_), .B(_17045_), .C(_17048_), .Y(_16897__25_) );
NOR3X1 NOR3X1_507 ( .gnd(gnd), .vdd(vdd), .A(_16904_), .B(_16924_), .C(_17001_), .Y(_17049_) );
XNOR2X1 XNOR2X1_446 ( .gnd(gnd), .vdd(vdd), .A(_17049_), .B(module_3_W_26_), .Y(_17050_) );
NOR2X1 NOR2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf7), .B(nonce_iniciales[122]), .Y(_17051_) );
AOI21X1 AOI21X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_16933__bF_buf2), .B(_17050_), .C(_17051_), .Y(_16897__26_) );
NOR2X1 NOR2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[123]), .Y(_17052_) );
AND2X2 AND2X2_387 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_26_), .B(module_3_W_25_), .Y(_17053_) );
NAND3X1 NAND3X1_3909 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_24_), .B(_17053_), .C(_17040_), .Y(_17054_) );
OR2X2 OR2X2_412 ( .gnd(gnd), .vdd(vdd), .A(_17054_), .B(module_3_W_27_), .Y(_17055_) );
AOI21X1 AOI21X1_2426 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_27_), .B(_17054_), .C(_16970_), .Y(_17056_) );
AOI21X1 AOI21X1_2427 ( .gnd(gnd), .vdd(vdd), .A(_17055_), .B(_17056_), .C(_17052_), .Y(_16897__27_) );
INVX1 INVX1_2414 ( .gnd(gnd), .vdd(vdd), .A(_16906_), .Y(_17057_) );
NOR3X1 NOR3X1_508 ( .gnd(gnd), .vdd(vdd), .A(_17057_), .B(_16924_), .C(_17001_), .Y(_17058_) );
NAND2X1 NAND2X1_2269 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_28_), .B(_17058_), .Y(_17059_) );
INVX1 INVX1_2415 ( .gnd(gnd), .vdd(vdd), .A(_16924_), .Y(_17060_) );
NAND3X1 NAND3X1_3910 ( .gnd(gnd), .vdd(vdd), .A(_16906_), .B(_17060_), .C(_16995_), .Y(_17061_) );
NAND2X1 NAND2X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_16911_), .B(_17061_), .Y(_17062_) );
NAND2X1 NAND2X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_17059_), .B(_17062_), .Y(_17063_) );
NOR2X1 NOR2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf6), .B(nonce_iniciales[124]), .Y(_17064_) );
AOI21X1 AOI21X1_2428 ( .gnd(gnd), .vdd(vdd), .A(_16933__bF_buf0), .B(_17063_), .C(_17064_), .Y(_16897__28_) );
NOR2X1 NOR2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf6), .B(nonce_iniciales[125]), .Y(_17065_) );
OR2X2 OR2X2_413 ( .gnd(gnd), .vdd(vdd), .A(_17059_), .B(module_3_W_29_), .Y(_17066_) );
AOI21X1 AOI21X1_2429 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_29_), .B(_17059_), .C(_16970_), .Y(_17067_) );
AOI21X1 AOI21X1_2430 ( .gnd(gnd), .vdd(vdd), .A(_17066_), .B(_17067_), .C(_17065_), .Y(_16897__29_) );
NAND3X1 NAND3X1_3911 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_30_), .B(_16912_), .C(_17058_), .Y(_17068_) );
INVX1 INVX1_2416 ( .gnd(gnd), .vdd(vdd), .A(_16912_), .Y(_17069_) );
OAI21X1 OAI21X1_2741 ( .gnd(gnd), .vdd(vdd), .A(_17061_), .B(_17069_), .C(_16914_), .Y(_17070_) );
NAND2X1 NAND2X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_17068_), .B(_17070_), .Y(_17071_) );
NOR2X1 NOR2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[126]), .Y(_17072_) );
AOI21X1 AOI21X1_2431 ( .gnd(gnd), .vdd(vdd), .A(_16933__bF_buf0), .B(_17071_), .C(_17072_), .Y(_16897__30_) );
NOR2X1 NOR2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(inicio_bF_buf4), .B(nonce_iniciales[127]), .Y(_17073_) );
NOR2X1 NOR2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_17069_), .B(_17061_), .Y(_17074_) );
NAND3X1 NAND3X1_3912 ( .gnd(gnd), .vdd(vdd), .A(_16913_), .B(module_3_W_30_), .C(_17074_), .Y(_17075_) );
AOI21X1 AOI21X1_2432 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_31_), .B(_17068_), .C(_16970_), .Y(_17076_) );
AOI21X1 AOI21X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_17075_), .B(_17076_), .C(_17073_), .Y(_16897__31_) );
DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_16897__0_), .Q(module_3_W_0_) );
DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_16897__1_), .Q(module_3_W_1_) );
DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_16897__2_), .Q(module_3_W_2_) );
DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_16897__3_), .Q(module_3_W_3_) );
DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_16897__4_), .Q(module_3_W_4_) );
DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_16897__5_), .Q(module_3_W_5_) );
DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_16897__6_), .Q(module_3_W_6_) );
DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_16897__7_), .Q(module_3_W_7_) );
DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_16897__8_), .Q(module_3_W_8_) );
DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_16897__9_), .Q(module_3_W_9_) );
DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_16897__10_), .Q(module_3_W_10_) );
DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_16897__11_), .Q(module_3_W_11_) );
DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__12_), .Q(module_3_W_12_) );
DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_16897__13_), .Q(module_3_W_13_) );
DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__14_), .Q(module_3_W_14_) );
DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__15_), .Q(module_3_W_15_) );
DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_16897__16_), .Q(module_3_W_16_) );
DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__17_), .Q(module_3_W_17_) );
DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__18_), .Q(module_3_W_18_) );
DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__19_), .Q(module_3_W_19_) );
DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_16897__20_), .Q(module_3_W_20_) );
DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__21_), .Q(module_3_W_21_) );
DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__22_), .Q(module_3_W_22_) );
DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__23_), .Q(module_3_W_23_) );
DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_16897__24_), .Q(module_3_W_24_) );
DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__25_), .Q(module_3_W_25_) );
DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__26_), .Q(module_3_W_26_) );
DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_16897__27_), .Q(module_3_W_27_) );
DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_16897__28_), .Q(module_3_W_28_) );
DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_16897__29_), .Q(module_3_W_29_) );
DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_16897__30_), .Q(module_3_W_30_) );
DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_16897__31_), .Q(module_3_W_31_) );
INVX1 INVX1_2417 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_17116_) );
INVX1 INVX1_2418 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .Y(_17117_) );
INVX1 INVX1_2419 ( .gnd(gnd), .vdd(vdd), .A(target[0]), .Y(_17118_) );
OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_17117_), .B(gnd), .C(_17118_), .D(vdd), .Y(_17119_) );
OAI21X1 OAI21X1_2742 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .B(_17116_), .C(_17119_), .Y(_17120_) );
XOR2X1 XOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(vdd), .Y(_17121_) );
INVX2 INVX2_602 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .Y(_17122_) );
INVX1 INVX1_2420 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_17123_) );
NAND2X1 NAND2X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_17122_), .B(_17123_), .Y(_17124_) );
NAND2X1 NAND2X1_2274 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(gnd), .Y(_17125_) );
AOI21X1 AOI21X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_17124_), .B(_17125_), .C(_17121_), .Y(_17126_) );
INVX1 INVX1_2421 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .Y(_17127_) );
NAND2X1 NAND2X1_2275 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(_17127_), .Y(_17128_) );
NAND2X1 NAND2X1_2276 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_17122_), .Y(_17129_) );
OAI21X1 OAI21X1_2743 ( .gnd(gnd), .vdd(vdd), .A(_17121_), .B(_17129_), .C(_17128_), .Y(_17130_) );
AOI21X1 AOI21X1_2435 ( .gnd(gnd), .vdd(vdd), .A(_17120_), .B(_17126_), .C(_17130_), .Y(_17131_) );
INVX1 INVX1_2422 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_15_), .Y(_17132_) );
INVX1 INVX1_2423 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_14_), .Y(_17133_) );
OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_17132_), .B(target[7]), .C(target[6]), .D(_17133_), .Y(_17134_) );
INVX4 INVX4_16 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .Y(_17135_) );
INVX2 INVX2_603 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .Y(_17136_) );
OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_17135_), .B(module_3_H_15_), .C(_17136_), .D(module_3_H_14_), .Y(_17137_) );
NOR2X1 NOR2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_17134_), .B(_17137_), .Y(_17138_) );
INVX2 INVX2_604 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_13_), .Y(_17139_) );
INVX1 INVX1_2424 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_12_), .Y(_17140_) );
OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_17139_), .B(target[5]), .C(target[4]), .D(_17140_), .Y(_17141_) );
INVX2 INVX2_605 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .Y(_17142_) );
INVX1 INVX1_2425 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .Y(_17143_) );
OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_17142_), .B(module_3_H_13_), .C(_17143_), .D(module_3_H_12_), .Y(_17144_) );
NOR2X1 NOR2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_17141_), .B(_17144_), .Y(_17145_) );
NAND2X1 NAND2X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_17138_), .B(_17145_), .Y(_17146_) );
NAND2X1 NAND2X1_2278 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .B(_17139_), .Y(_17147_) );
NAND3X1 NAND3X1_3913 ( .gnd(gnd), .vdd(vdd), .A(_17141_), .B(_17147_), .C(_17138_), .Y(_17148_) );
OAI21X1 OAI21X1_2744 ( .gnd(gnd), .vdd(vdd), .A(_17131_), .B(_17146_), .C(_17148_), .Y(_17149_) );
INVX1 INVX1_2426 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_17_), .Y(_17150_) );
OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_17117_), .B(module_3_H_17_), .C(_17118_), .D(module_3_H_16_), .Y(_17151_) );
OAI21X1 OAI21X1_2745 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .B(_17150_), .C(_17151_), .Y(_17152_) );
XOR2X1 XOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(module_3_H_19_), .Y(_17153_) );
INVX1 INVX1_2427 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_18_), .Y(_17154_) );
NAND2X1 NAND2X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_17122_), .B(_17154_), .Y(_17155_) );
NAND2X1 NAND2X1_2280 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(module_3_H_18_), .Y(_17156_) );
AOI21X1 AOI21X1_2436 ( .gnd(gnd), .vdd(vdd), .A(_17155_), .B(_17156_), .C(_17153_), .Y(_17157_) );
NAND2X1 NAND2X1_2281 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_19_), .B(_17127_), .Y(_17079_) );
NAND2X1 NAND2X1_2282 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_18_), .B(_17122_), .Y(_17080_) );
OAI21X1 OAI21X1_2746 ( .gnd(gnd), .vdd(vdd), .A(_17153_), .B(_17080_), .C(_17079_), .Y(_17081_) );
AOI21X1 AOI21X1_2437 ( .gnd(gnd), .vdd(vdd), .A(_17152_), .B(_17157_), .C(_17081_), .Y(_17082_) );
INVX1 INVX1_2428 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_23_), .Y(_17083_) );
INVX1 INVX1_2429 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_22_), .Y(_17084_) );
OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_17083_), .B(target[7]), .C(target[6]), .D(_17084_), .Y(_17085_) );
OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_17135_), .B(module_3_H_23_), .C(_17136_), .D(module_3_H_22_), .Y(_17086_) );
NOR2X1 NOR2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_17085_), .B(_17086_), .Y(_17087_) );
NAND2X1 NAND2X1_2283 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_21_), .B(_17142_), .Y(_17088_) );
NAND2X1 NAND2X1_2284 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_20_), .B(_17143_), .Y(_17089_) );
AND2X2 AND2X2_388 ( .gnd(gnd), .vdd(vdd), .A(_17088_), .B(_17089_), .Y(_17090_) );
INVX1 INVX1_2430 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_20_), .Y(_17091_) );
NOR2X1 NOR2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_21_), .B(_17142_), .Y(_17092_) );
AOI21X1 AOI21X1_2438 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_17091_), .C(_17092_), .Y(_17093_) );
NAND3X1 NAND3X1_3914 ( .gnd(gnd), .vdd(vdd), .A(_17090_), .B(_17093_), .C(_17087_), .Y(_17094_) );
AOI21X1 AOI21X1_2439 ( .gnd(gnd), .vdd(vdd), .A(_17088_), .B(_17089_), .C(_17092_), .Y(_17095_) );
AOI22X1 AOI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_17135_), .B(module_3_H_23_), .C(_17136_), .D(module_3_H_22_), .Y(_17096_) );
NOR2X1 NOR2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_23_), .B(_17135_), .Y(_17097_) );
AOI22X1 AOI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_17135_), .B(module_3_H_15_), .C(_17136_), .D(module_3_H_14_), .Y(_17098_) );
NOR2X1 NOR2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_15_), .B(_17135_), .Y(_17099_) );
OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_17096_), .B(_17097_), .C(_17098_), .D(_17099_), .Y(_17100_) );
AOI21X1 AOI21X1_2440 ( .gnd(gnd), .vdd(vdd), .A(_17087_), .B(_17095_), .C(_17100_), .Y(_17101_) );
OAI21X1 OAI21X1_2747 ( .gnd(gnd), .vdd(vdd), .A(_17082_), .B(_17094_), .C(_17101_), .Y(_17102_) );
NOR2X1 NOR2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf2), .B(_17102__bF_buf3), .Y(module_3_comparador_target_hash_0_terminado) );
INVX1 INVX1_2431 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_0_), .Y(_17103_) );
NOR3X1 NOR3X1_509 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf2), .B(_17103_), .C(_17102__bF_buf3), .Y(bounty_72_) );
INVX1 INVX1_2432 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_1_), .Y(_17104_) );
NOR3X1 NOR3X1_510 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf1), .B(_17104_), .C(_17102__bF_buf0), .Y(bounty_73_) );
INVX1 INVX1_2433 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_2_), .Y(_17105_) );
NOR3X1 NOR3X1_511 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf1), .B(_17105_), .C(_17102__bF_buf0), .Y(bounty_74_) );
INVX1 INVX1_2434 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_3_), .Y(_17106_) );
NOR3X1 NOR3X1_512 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf1), .B(_17106_), .C(_17102__bF_buf0), .Y(bounty_75_) );
INVX1 INVX1_2435 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_4_), .Y(_17107_) );
NOR3X1 NOR3X1_513 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf2), .B(_17107_), .C(_17102__bF_buf3), .Y(bounty_76_) );
INVX1 INVX1_2436 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_5_), .Y(_17108_) );
NOR3X1 NOR3X1_514 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf1), .B(_17108_), .C(_17102__bF_buf0), .Y(bounty_77_) );
INVX1 INVX1_2437 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_6_), .Y(_17109_) );
NOR3X1 NOR3X1_515 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf0), .B(_17109_), .C(_17102__bF_buf1), .Y(bounty_78_) );
INVX1 INVX1_2438 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_7_), .Y(_17110_) );
NOR3X1 NOR3X1_516 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf3), .B(_17110_), .C(_17102__bF_buf4), .Y(bounty_79_) );
INVX1 INVX1_2439 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_17111_) );
NOR3X1 NOR3X1_517 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf3), .B(_17111_), .C(_17102__bF_buf4), .Y(bounty_80_) );
NOR3X1 NOR3X1_518 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf3), .B(_17116_), .C(_17102__bF_buf4), .Y(bounty_81_) );
NOR3X1 NOR3X1_519 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf4), .B(_17123_), .C(_17102__bF_buf2), .Y(bounty_82_) );
INVX1 INVX1_2440 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_17112_) );
NOR3X1 NOR3X1_520 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf4), .B(_17112_), .C(_17102__bF_buf1), .Y(bounty_83_) );
NOR3X1 NOR3X1_521 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf3), .B(_17140_), .C(_17102__bF_buf4), .Y(bounty_84_) );
NOR3X1 NOR3X1_522 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf2), .B(_17139_), .C(_17102__bF_buf3), .Y(bounty_85_) );
NOR3X1 NOR3X1_523 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf1), .B(_17133_), .C(_17102__bF_buf0), .Y(bounty_86_) );
NOR3X1 NOR3X1_524 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf2), .B(_17132_), .C(_17102__bF_buf3), .Y(bounty_87_) );
INVX1 INVX1_2441 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_16_), .Y(_17113_) );
NOR3X1 NOR3X1_525 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf4), .B(_17113_), .C(_17102__bF_buf2), .Y(bounty_88_) );
NOR3X1 NOR3X1_526 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf0), .B(_17150_), .C(_17102__bF_buf2), .Y(bounty_89_) );
NOR3X1 NOR3X1_527 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf4), .B(_17154_), .C(_17102__bF_buf2), .Y(bounty_90_) );
INVX1 INVX1_2442 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_19_), .Y(_17114_) );
NOR3X1 NOR3X1_528 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf4), .B(_17114_), .C(_17102__bF_buf2), .Y(bounty_91_) );
NOR3X1 NOR3X1_529 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf0), .B(_17091_), .C(_17102__bF_buf1), .Y(bounty_92_) );
INVX1 INVX1_2443 ( .gnd(gnd), .vdd(vdd), .A(module_3_H_21_), .Y(_17115_) );
NOR3X1 NOR3X1_530 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf3), .B(_17115_), .C(_17102__bF_buf4), .Y(bounty_93_) );
NOR3X1 NOR3X1_531 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf0), .B(_17084_), .C(_17102__bF_buf1), .Y(bounty_94_) );
NOR3X1 NOR3X1_532 ( .gnd(gnd), .vdd(vdd), .A(_17149__bF_buf0), .B(_17083_), .C(_17102__bF_buf1), .Y(bounty_95_) );
INVX1 INVX1_2444 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf3_), .Y(_17158_) );
AOI21X1 AOI21X1_2441 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_24_), .B(_17158_), .C(bloque_datos_80_bF_buf2_), .Y(_17159_) );
OAI21X1 OAI21X1_2748 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_24_), .B(_17158_), .C(_17159_), .Y(module_3_W_136_) );
INVX1 INVX1_2445 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf3_), .Y(_17160_) );
AOI21X1 AOI21X1_2442 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_25_), .B(_17160_), .C(bloque_datos_81_bF_buf4_), .Y(_17161_) );
OAI21X1 OAI21X1_2749 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_25_), .B(_17160_), .C(_17161_), .Y(module_3_W_137_) );
INVX1 INVX1_2446 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf3_), .Y(_17162_) );
AOI21X1 AOI21X1_2443 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_26_), .B(_17162_), .C(bloque_datos_82_bF_buf1_), .Y(_17163_) );
OAI21X1 OAI21X1_2750 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_26_), .B(_17162_), .C(_17163_), .Y(module_3_W_138_) );
INVX1 INVX1_2447 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf3_), .Y(_17164_) );
AOI21X1 AOI21X1_2444 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_27_), .B(_17164_), .C(bloque_datos_83_bF_buf2_), .Y(_17165_) );
OAI21X1 OAI21X1_2751 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_27_), .B(_17164_), .C(_17165_), .Y(module_3_W_139_) );
INVX1 INVX1_2448 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf1_), .Y(_17166_) );
AOI21X1 AOI21X1_2445 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_28_), .B(_17166_), .C(bloque_datos_84_bF_buf3_), .Y(_17167_) );
OAI21X1 OAI21X1_2752 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_28_), .B(_17166_), .C(_17167_), .Y(module_3_W_140_) );
INVX1 INVX1_2449 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf1_), .Y(_17168_) );
AOI21X1 AOI21X1_2446 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_29_), .B(_17168_), .C(bloque_datos_85_bF_buf0_), .Y(_17169_) );
OAI21X1 OAI21X1_2753 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_29_), .B(_17168_), .C(_17169_), .Y(module_3_W_141_) );
INVX1 INVX1_2450 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf1_), .Y(_17170_) );
AOI21X1 AOI21X1_2447 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_30_), .B(_17170_), .C(bloque_datos_86_bF_buf3_), .Y(_17171_) );
OAI21X1 OAI21X1_2754 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_30_), .B(_17170_), .C(_17171_), .Y(module_3_W_142_) );
INVX1 INVX1_2451 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .Y(_17172_) );
AOI21X1 AOI21X1_2448 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_31_), .B(_17172_), .C(bloque_datos_87_bF_buf2_), .Y(_17173_) );
OAI21X1 OAI21X1_2755 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_31_), .B(_17172_), .C(_17173_), .Y(module_3_W_143_) );
INVX1 INVX1_2452 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf4_), .Y(_17174_) );
OR2X2 OR2X2_414 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_16_), .B(bloque_datos_24_bF_buf3_), .Y(_17175_) );
NAND2X1 NAND2X1_2285 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_16_), .B(bloque_datos_24_bF_buf2_), .Y(_17176_) );
NAND2X1 NAND2X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_17176_), .B(_17175_), .Y(_17177_) );
NAND2X1 NAND2X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_17174_), .B(_17177_), .Y(module_3_W_128_) );
INVX1 INVX1_2453 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf2_), .Y(_17178_) );
AOI21X1 AOI21X1_2449 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_17_), .B(_17178_), .C(bloque_datos_73_bF_buf2_), .Y(_17179_) );
OAI21X1 OAI21X1_2756 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_17_), .B(_17178_), .C(_17179_), .Y(module_3_W_129_) );
INVX1 INVX1_2454 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf4_), .Y(_17180_) );
OR2X2 OR2X2_415 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_18_), .B(bloque_datos_26_bF_buf2_), .Y(_17181_) );
NAND2X1 NAND2X1_2288 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_18_), .B(bloque_datos_26_bF_buf1_), .Y(_17182_) );
NAND2X1 NAND2X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_17182_), .B(_17181_), .Y(_17183_) );
NAND2X1 NAND2X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_17180_), .B(_17183_), .Y(module_3_W_130_) );
INVX1 INVX1_2455 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf0_), .Y(_17184_) );
OR2X2 OR2X2_416 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_19_), .B(bloque_datos_27_bF_buf0_), .Y(_17185_) );
NAND2X1 NAND2X1_2291 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_19_), .B(bloque_datos_27_bF_buf4_), .Y(_17186_) );
NAND2X1 NAND2X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_17186_), .B(_17185_), .Y(_17187_) );
NAND2X1 NAND2X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_17184_), .B(_17187_), .Y(module_3_W_131_) );
INVX2 INVX2_606 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf0_), .Y(_17188_) );
AOI21X1 AOI21X1_2450 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_20_), .B(_17188_), .C(bloque_datos_76_bF_buf3_), .Y(_17189_) );
OAI21X1 OAI21X1_2757 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_20_), .B(_17188_), .C(_17189_), .Y(module_3_W_132_) );
INVX2 INVX2_607 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf0_), .Y(_17190_) );
AOI21X1 AOI21X1_2451 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_21_), .B(_17190_), .C(bloque_datos_77_bF_buf3_), .Y(_17191_) );
OAI21X1 OAI21X1_2758 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_21_), .B(_17190_), .C(_17191_), .Y(module_3_W_133_) );
INVX2 INVX2_608 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf1_), .Y(_17192_) );
AOI21X1 AOI21X1_2452 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_22_), .B(_17192_), .C(bloque_datos_78_bF_buf3_), .Y(_17193_) );
OAI21X1 OAI21X1_2759 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_22_), .B(_17192_), .C(_17193_), .Y(module_3_W_134_) );
INVX1 INVX1_2456 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf1_), .Y(_17194_) );
AOI21X1 AOI21X1_2453 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_23_), .B(_17194_), .C(bloque_datos_79_bF_buf2_), .Y(_17195_) );
OAI21X1 OAI21X1_2760 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_23_), .B(_17194_), .C(_17195_), .Y(module_3_W_135_) );
INVX1 INVX1_2457 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(_17196_) );
INVX1 INVX1_2458 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf0_), .Y(_17197_) );
OAI21X1 OAI21X1_2761 ( .gnd(gnd), .vdd(vdd), .A(_17196_), .B(bloque_datos_40_bF_buf3_), .C(_17197_), .Y(_17198_) );
AOI21X1 AOI21X1_2454 ( .gnd(gnd), .vdd(vdd), .A(_17196_), .B(bloque_datos_40_bF_buf2_), .C(_17198_), .Y(_17199_) );
INVX1 INVX1_2459 ( .gnd(gnd), .vdd(vdd), .A(_17199_), .Y(module_3_W_144_) );
INVX1 INVX1_2460 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(_17200_) );
INVX1 INVX1_2461 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf3_), .Y(_17201_) );
OAI21X1 OAI21X1_2762 ( .gnd(gnd), .vdd(vdd), .A(_17200_), .B(bloque_datos_41_bF_buf2_), .C(_17201_), .Y(_17202_) );
AOI21X1 AOI21X1_2455 ( .gnd(gnd), .vdd(vdd), .A(_17200_), .B(bloque_datos_41_bF_buf1_), .C(_17202_), .Y(_17203_) );
INVX1 INVX1_2462 ( .gnd(gnd), .vdd(vdd), .A(_17203_), .Y(module_3_W_145_) );
INVX1 INVX1_2463 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf0_), .Y(_17204_) );
INVX1 INVX1_2464 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf0_), .Y(_17205_) );
OAI21X1 OAI21X1_2763 ( .gnd(gnd), .vdd(vdd), .A(_17204_), .B(bloque_datos_42_bF_buf2_), .C(_17205_), .Y(_17206_) );
AOI21X1 AOI21X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_17204_), .B(bloque_datos_42_bF_buf1_), .C(_17206_), .Y(_17207_) );
INVX1 INVX1_2465 ( .gnd(gnd), .vdd(vdd), .A(_17207_), .Y(module_3_W_146_) );
INVX1 INVX1_2466 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf0_), .Y(_17208_) );
INVX1 INVX1_2467 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf1_), .Y(_17209_) );
OAI21X1 OAI21X1_2764 ( .gnd(gnd), .vdd(vdd), .A(_17208_), .B(bloque_datos_43_bF_buf2_), .C(_17209_), .Y(_17210_) );
AOI21X1 AOI21X1_2457 ( .gnd(gnd), .vdd(vdd), .A(_17208_), .B(bloque_datos_43_bF_buf1_), .C(_17210_), .Y(_17211_) );
INVX1 INVX1_2468 ( .gnd(gnd), .vdd(vdd), .A(_17211_), .Y(module_3_W_147_) );
INVX1 INVX1_2469 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf0_), .Y(_17212_) );
INVX1 INVX1_2470 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf0_), .Y(_17213_) );
OAI21X1 OAI21X1_2765 ( .gnd(gnd), .vdd(vdd), .A(_17212_), .B(bloque_datos_44_bF_buf3_), .C(_17213_), .Y(_17214_) );
AOI21X1 AOI21X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_17212_), .B(bloque_datos_44_bF_buf2_), .C(_17214_), .Y(_17215_) );
INVX1 INVX1_2471 ( .gnd(gnd), .vdd(vdd), .A(_17215_), .Y(module_3_W_148_) );
INVX1 INVX1_2472 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf0_), .Y(_17216_) );
INVX1 INVX1_2473 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf0_), .Y(_17217_) );
OAI21X1 OAI21X1_2766 ( .gnd(gnd), .vdd(vdd), .A(_17216_), .B(bloque_datos_45_bF_buf3_), .C(_17217_), .Y(_17218_) );
AOI21X1 AOI21X1_2459 ( .gnd(gnd), .vdd(vdd), .A(_17216_), .B(bloque_datos_45_bF_buf2_), .C(_17218_), .Y(_17219_) );
INVX1 INVX1_2474 ( .gnd(gnd), .vdd(vdd), .A(_17219_), .Y(module_3_W_149_) );
INVX1 INVX1_2475 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf0_), .Y(_17220_) );
INVX1 INVX1_2476 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf0_), .Y(_17221_) );
OAI21X1 OAI21X1_2767 ( .gnd(gnd), .vdd(vdd), .A(_17220_), .B(bloque_datos_46_bF_buf3_), .C(_17221_), .Y(_17222_) );
AOI21X1 AOI21X1_2460 ( .gnd(gnd), .vdd(vdd), .A(_17220_), .B(bloque_datos_46_bF_buf2_), .C(_17222_), .Y(_17223_) );
INVX2 INVX2_609 ( .gnd(gnd), .vdd(vdd), .A(_17223_), .Y(module_3_W_150_) );
INVX1 INVX1_2477 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[7]), .Y(_17224_) );
INVX1 INVX1_2478 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf1_), .Y(_17225_) );
OAI21X1 OAI21X1_2768 ( .gnd(gnd), .vdd(vdd), .A(_17224_), .B(bloque_datos_47_bF_buf2_), .C(_17225_), .Y(_17226_) );
AOI21X1 AOI21X1_2461 ( .gnd(gnd), .vdd(vdd), .A(_17224_), .B(bloque_datos_47_bF_buf1_), .C(_17226_), .Y(_17227_) );
INVX2 INVX2_610 ( .gnd(gnd), .vdd(vdd), .A(_17227_), .Y(module_3_W_151_) );
AOI21X1 AOI21X1_2462 ( .gnd(gnd), .vdd(vdd), .A(_17176_), .B(_17175_), .C(bloque_datos_72_bF_buf3_), .Y(_17228_) );
XNOR2X1 XNOR2X1_447 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .B(bloque_datos_48_bF_buf3_), .Y(_17229_) );
NAND2X1 NAND2X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_17229_), .B(_17228_), .Y(module_3_W_152_) );
XOR2X1 XOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .B(bloque_datos_49_bF_buf2_), .Y(_17230_) );
NOR2X1 NOR2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_17230_), .B(module_3_W_129_), .Y(_17231_) );
INVX1 INVX1_2479 ( .gnd(gnd), .vdd(vdd), .A(_17231_), .Y(module_3_W_153_) );
AOI21X1 AOI21X1_2463 ( .gnd(gnd), .vdd(vdd), .A(_17182_), .B(_17181_), .C(bloque_datos_74_bF_buf3_), .Y(_17232_) );
XNOR2X1 XNOR2X1_448 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .B(bloque_datos_50_bF_buf2_), .Y(_17233_) );
NAND2X1 NAND2X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_17233_), .B(_17232_), .Y(module_3_W_154_) );
AOI21X1 AOI21X1_2464 ( .gnd(gnd), .vdd(vdd), .A(_17186_), .B(_17185_), .C(bloque_datos_75_bF_buf4_), .Y(_17234_) );
XNOR2X1 XNOR2X1_449 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .B(bloque_datos_51_bF_buf2_), .Y(_17235_) );
NAND2X1 NAND2X1_2296 ( .gnd(gnd), .vdd(vdd), .A(_17235_), .B(_17234_), .Y(module_3_W_155_) );
INVX1 INVX1_2480 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_20_), .Y(_17236_) );
INVX1 INVX1_2481 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf2_), .Y(_17237_) );
OAI21X1 OAI21X1_2769 ( .gnd(gnd), .vdd(vdd), .A(_17236_), .B(bloque_datos_28_bF_buf4_), .C(_17237_), .Y(_17238_) );
AOI21X1 AOI21X1_2465 ( .gnd(gnd), .vdd(vdd), .A(_17236_), .B(bloque_datos_28_bF_buf3_), .C(_17238_), .Y(_17239_) );
AND2X2 AND2X2_389 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf1_), .B(bloque_datos_52_bF_buf3_), .Y(_17240_) );
NOR2X1 NOR2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf0_), .B(bloque_datos_52_bF_buf2_), .Y(_17241_) );
OAI21X1 OAI21X1_2770 ( .gnd(gnd), .vdd(vdd), .A(_17240_), .B(_17241_), .C(_17239_), .Y(module_3_W_156_) );
XOR2X1 XOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf0_), .B(bloque_datos_53_bF_buf1_), .Y(_17242_) );
NOR2X1 NOR2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_17242_), .B(module_3_W_133_), .Y(_17243_) );
INVX1 INVX1_2482 ( .gnd(gnd), .vdd(vdd), .A(_17243_), .Y(module_3_W_157_) );
XOR2X1 XOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf0_), .B(bloque_datos_54_bF_buf1_), .Y(_17244_) );
NOR2X1 NOR2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_17244_), .B(module_3_W_134_), .Y(_17245_) );
INVX1 INVX1_2483 ( .gnd(gnd), .vdd(vdd), .A(_17245_), .Y(module_3_W_158_) );
XOR2X1 XOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[15]), .B(bloque_datos[55]), .Y(_17246_) );
NOR2X1 NOR2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_17246_), .B(module_3_W_135_), .Y(_17247_) );
INVX1 INVX1_2484 ( .gnd(gnd), .vdd(vdd), .A(_17247_), .Y(module_3_W_159_) );
XOR2X1 XOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_24_), .B(bloque_datos_32_bF_buf2_), .Y(_17248_) );
NOR2X1 NOR2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf1_), .B(_17248_), .Y(_17249_) );
XNOR2X1 XNOR2X1_450 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf0_), .B(bloque_datos_56_bF_buf3_), .Y(_17250_) );
NAND2X1 NAND2X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_17250_), .B(_17249_), .Y(module_3_W_160_) );
INVX1 INVX1_2485 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_25_), .Y(_17251_) );
INVX1 INVX1_2486 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf3_), .Y(_17252_) );
OAI21X1 OAI21X1_2771 ( .gnd(gnd), .vdd(vdd), .A(_17251_), .B(bloque_datos_33_bF_buf2_), .C(_17252_), .Y(_17253_) );
AOI21X1 AOI21X1_2466 ( .gnd(gnd), .vdd(vdd), .A(_17251_), .B(bloque_datos_33_bF_buf1_), .C(_17253_), .Y(_17254_) );
XNOR2X1 XNOR2X1_451 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .B(bloque_datos_57_bF_buf2_), .Y(_17255_) );
NAND2X1 NAND2X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_17255_), .B(_17254_), .Y(module_3_W_161_) );
XOR2X1 XOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_26_), .B(bloque_datos_34_bF_buf2_), .Y(_17256_) );
NOR2X1 NOR2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf0_), .B(_17256_), .Y(_17257_) );
XNOR2X1 XNOR2X1_452 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .B(bloque_datos_58_bF_buf3_), .Y(_17258_) );
NAND2X1 NAND2X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_17258_), .B(_17257_), .Y(module_3_W_162_) );
XOR2X1 XOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_27_), .B(bloque_datos_35_bF_buf2_), .Y(_17259_) );
NOR2X1 NOR2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf1_), .B(_17259_), .Y(_17260_) );
XNOR2X1 XNOR2X1_453 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf0_), .B(bloque_datos_59_bF_buf3_), .Y(_17261_) );
NAND2X1 NAND2X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_17261_), .B(_17260_), .Y(module_3_W_163_) );
XOR2X1 XOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf0_), .B(bloque_datos_60_bF_buf1_), .Y(_17262_) );
NOR2X1 NOR2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_17262_), .B(module_3_W_140_), .Y(_17263_) );
INVX1 INVX1_2487 ( .gnd(gnd), .vdd(vdd), .A(_17263_), .Y(module_3_W_164_) );
XOR2X1 XOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf0_), .B(bloque_datos_61_bF_buf3_), .Y(_17264_) );
NOR2X1 NOR2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_17264_), .B(module_3_W_141_), .Y(_17265_) );
INVX1 INVX1_2488 ( .gnd(gnd), .vdd(vdd), .A(_17265_), .Y(module_3_W_165_) );
XOR2X1 XOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf0_), .B(bloque_datos_62_bF_buf1_), .Y(_17266_) );
NOR2X1 NOR2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_17266_), .B(module_3_W_142_), .Y(_17267_) );
INVX2 INVX2_611 ( .gnd(gnd), .vdd(vdd), .A(_17267_), .Y(module_3_W_166_) );
XOR2X1 XOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf0_), .B(bloque_datos[63]), .Y(_17268_) );
NOR2X1 NOR2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_17268_), .B(module_3_W_143_), .Y(_17269_) );
INVX1 INVX1_2489 ( .gnd(gnd), .vdd(vdd), .A(_17269_), .Y(module_3_W_167_) );
XNOR2X1 XNOR2X1_454 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf1_), .B(bloque_datos_64_bF_buf3_), .Y(_17270_) );
AND2X2 AND2X2_390 ( .gnd(gnd), .vdd(vdd), .A(_17199_), .B(_17270_), .Y(_17271_) );
INVX2 INVX2_612 ( .gnd(gnd), .vdd(vdd), .A(_17271_), .Y(module_3_W_168_) );
XNOR2X1 XNOR2X1_455 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf1_), .B(bloque_datos_65_bF_buf2_), .Y(_17272_) );
AND2X2 AND2X2_391 ( .gnd(gnd), .vdd(vdd), .A(_17203_), .B(_17272_), .Y(_17273_) );
INVX1 INVX1_2490 ( .gnd(gnd), .vdd(vdd), .A(_17273_), .Y(module_3_W_169_) );
XNOR2X1 XNOR2X1_456 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf0_), .B(bloque_datos_66_bF_buf3_), .Y(_17274_) );
AND2X2 AND2X2_392 ( .gnd(gnd), .vdd(vdd), .A(_17207_), .B(_17274_), .Y(_17275_) );
INVX1 INVX1_2491 ( .gnd(gnd), .vdd(vdd), .A(_17275_), .Y(module_3_W_170_) );
AND2X2 AND2X2_393 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf3_), .B(bloque_datos_67_bF_buf0_), .Y(_17276_) );
NOR2X1 NOR2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf2_), .B(bloque_datos_67_bF_buf4_), .Y(_17277_) );
OAI21X1 OAI21X1_2772 ( .gnd(gnd), .vdd(vdd), .A(_17276_), .B(_17277_), .C(_17211_), .Y(module_3_W_171_) );
INVX2 INVX2_613 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf1_), .Y(_17278_) );
NOR2X1 NOR2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_17188_), .B(_17278_), .Y(_17279_) );
NOR2X1 NOR2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf2_), .B(bloque_datos_68_bF_buf0_), .Y(_17280_) );
OAI21X1 OAI21X1_2773 ( .gnd(gnd), .vdd(vdd), .A(_17279_), .B(_17280_), .C(_17215_), .Y(module_3_W_172_) );
INVX2 INVX2_614 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf1_), .Y(_17281_) );
NOR2X1 NOR2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_17190_), .B(_17281_), .Y(_17282_) );
NOR2X1 NOR2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf4_), .B(bloque_datos_69_bF_buf0_), .Y(_17283_) );
OAI21X1 OAI21X1_2774 ( .gnd(gnd), .vdd(vdd), .A(_17282_), .B(_17283_), .C(_17219_), .Y(module_3_W_173_) );
INVX2 INVX2_615 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf1_), .Y(_17284_) );
NOR2X1 NOR2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_17192_), .B(_17284_), .Y(_17285_) );
NOR2X1 NOR2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf0_), .B(bloque_datos_70_bF_buf0_), .Y(_17286_) );
OAI21X1 OAI21X1_2775 ( .gnd(gnd), .vdd(vdd), .A(_17285_), .B(_17286_), .C(_17223_), .Y(module_3_W_174_) );
XNOR2X1 XNOR2X1_457 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf0_), .B(bloque_datos_71_bF_buf1_), .Y(_17287_) );
AND2X2 AND2X2_394 ( .gnd(gnd), .vdd(vdd), .A(_17227_), .B(_17287_), .Y(_17288_) );
INVX1 INVX1_2492 ( .gnd(gnd), .vdd(vdd), .A(_17288_), .Y(module_3_W_175_) );
XNOR2X1 XNOR2X1_458 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf1_), .B(bloque_datos_72_bF_buf2_), .Y(_17289_) );
NAND3X1 NAND3X1_3915 ( .gnd(gnd), .vdd(vdd), .A(_17229_), .B(_17289_), .C(_17228_), .Y(module_3_W_176_) );
INVX1 INVX1_2493 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_17_), .Y(_17290_) );
NAND2X1 NAND2X1_2301 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf0_), .B(_17290_), .Y(_17291_) );
AND2X2 AND2X2_395 ( .gnd(gnd), .vdd(vdd), .A(_17179_), .B(_17291_), .Y(_17292_) );
INVX1 INVX1_2494 ( .gnd(gnd), .vdd(vdd), .A(_17230_), .Y(_17293_) );
XNOR2X1 XNOR2X1_459 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf0_), .B(bloque_datos_73_bF_buf1_), .Y(_17294_) );
NAND3X1 NAND3X1_3916 ( .gnd(gnd), .vdd(vdd), .A(_17293_), .B(_17294_), .C(_17292_), .Y(module_3_W_177_) );
XNOR2X1 XNOR2X1_460 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf1_), .B(bloque_datos_74_bF_buf2_), .Y(_17295_) );
NAND3X1 NAND3X1_3917 ( .gnd(gnd), .vdd(vdd), .A(_17233_), .B(_17295_), .C(_17232_), .Y(module_3_W_178_) );
XNOR2X1 XNOR2X1_461 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf1_), .B(bloque_datos_75_bF_buf3_), .Y(_17296_) );
NAND3X1 NAND3X1_3918 ( .gnd(gnd), .vdd(vdd), .A(_17235_), .B(_17296_), .C(_17234_), .Y(module_3_W_179_) );
XOR2X1 XOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf0_), .B(bloque_datos_76_bF_buf1_), .Y(_17297_) );
NOR2X1 NOR2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_17297_), .B(module_3_W_156_), .Y(_17298_) );
INVX1 INVX1_2495 ( .gnd(gnd), .vdd(vdd), .A(_17298_), .Y(module_3_W_180_) );
INVX1 INVX1_2496 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_21_), .Y(_17299_) );
INVX1 INVX1_2497 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf2_), .Y(_17300_) );
OAI21X1 OAI21X1_2776 ( .gnd(gnd), .vdd(vdd), .A(_17299_), .B(bloque_datos_29_bF_buf3_), .C(_17300_), .Y(_17301_) );
AOI21X1 AOI21X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_17299_), .B(bloque_datos_29_bF_buf2_), .C(_17301_), .Y(_17302_) );
INVX1 INVX1_2498 ( .gnd(gnd), .vdd(vdd), .A(_17242_), .Y(_17303_) );
XNOR2X1 XNOR2X1_462 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf0_), .B(bloque_datos_77_bF_buf1_), .Y(_17304_) );
NAND3X1 NAND3X1_3919 ( .gnd(gnd), .vdd(vdd), .A(_17303_), .B(_17304_), .C(_17302_), .Y(module_3_W_181_) );
XNOR2X1 XNOR2X1_463 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf0_), .B(bloque_datos_78_bF_buf2_), .Y(_17305_) );
AND2X2 AND2X2_396 ( .gnd(gnd), .vdd(vdd), .A(_17245_), .B(_17305_), .Y(_17306_) );
INVX2 INVX2_616 ( .gnd(gnd), .vdd(vdd), .A(_17306_), .Y(module_3_W_182_) );
XNOR2X1 XNOR2X1_464 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .B(bloque_datos_79_bF_buf1_), .Y(_17307_) );
AND2X2 AND2X2_397 ( .gnd(gnd), .vdd(vdd), .A(_17247_), .B(_17307_), .Y(_17308_) );
INVX2 INVX2_617 ( .gnd(gnd), .vdd(vdd), .A(_17308_), .Y(module_3_W_183_) );
XNOR2X1 XNOR2X1_465 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf0_), .B(bloque_datos_40_bF_buf1_), .Y(_17309_) );
NAND3X1 NAND3X1_3920 ( .gnd(gnd), .vdd(vdd), .A(_17250_), .B(_17309_), .C(_17249_), .Y(module_3_W_184_) );
XNOR2X1 XNOR2X1_466 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf2_), .B(bloque_datos_41_bF_buf0_), .Y(_17310_) );
NAND3X1 NAND3X1_3921 ( .gnd(gnd), .vdd(vdd), .A(_17255_), .B(_17310_), .C(_17254_), .Y(module_3_W_185_) );
XNOR2X1 XNOR2X1_467 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf4_), .B(bloque_datos_42_bF_buf0_), .Y(_17311_) );
NAND3X1 NAND3X1_3922 ( .gnd(gnd), .vdd(vdd), .A(_17258_), .B(_17311_), .C(_17257_), .Y(module_3_W_186_) );
XNOR2X1 XNOR2X1_468 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf0_), .B(bloque_datos_43_bF_buf0_), .Y(_17312_) );
NAND3X1 NAND3X1_3923 ( .gnd(gnd), .vdd(vdd), .A(_17261_), .B(_17312_), .C(_17260_), .Y(module_3_W_187_) );
XNOR2X1 XNOR2X1_469 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf2_), .B(bloque_datos_44_bF_buf1_), .Y(_17313_) );
AND2X2 AND2X2_398 ( .gnd(gnd), .vdd(vdd), .A(_17263_), .B(_17313_), .Y(_17314_) );
INVX1 INVX1_2499 ( .gnd(gnd), .vdd(vdd), .A(_17314_), .Y(module_3_W_188_) );
XNOR2X1 XNOR2X1_470 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf4_), .B(bloque_datos_45_bF_buf1_), .Y(_17315_) );
AND2X2 AND2X2_399 ( .gnd(gnd), .vdd(vdd), .A(_17265_), .B(_17315_), .Y(_17316_) );
INVX1 INVX1_2500 ( .gnd(gnd), .vdd(vdd), .A(_17316_), .Y(module_3_W_189_) );
XNOR2X1 XNOR2X1_471 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf2_), .B(bloque_datos_46_bF_buf1_), .Y(_17317_) );
AND2X2 AND2X2_400 ( .gnd(gnd), .vdd(vdd), .A(_17267_), .B(_17317_), .Y(_17318_) );
INVX1 INVX1_2501 ( .gnd(gnd), .vdd(vdd), .A(_17318_), .Y(module_3_W_190_) );
XNOR2X1 XNOR2X1_472 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf1_), .B(bloque_datos_47_bF_buf0_), .Y(_17319_) );
AND2X2 AND2X2_401 ( .gnd(gnd), .vdd(vdd), .A(_17269_), .B(_17319_), .Y(_17320_) );
INVX1 INVX1_2502 ( .gnd(gnd), .vdd(vdd), .A(_17320_), .Y(module_3_W_191_) );
AND2X2 AND2X2_402 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf4_), .B(bloque_datos_48_bF_buf2_), .Y(_17321_) );
NOR2X1 NOR2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf3_), .B(bloque_datos_48_bF_buf1_), .Y(_17322_) );
OAI21X1 OAI21X1_2777 ( .gnd(gnd), .vdd(vdd), .A(_17321_), .B(_17322_), .C(_17271_), .Y(module_3_W_192_) );
AND2X2 AND2X2_403 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf2_), .B(bloque_datos_49_bF_buf1_), .Y(_17323_) );
NOR2X1 NOR2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf1_), .B(bloque_datos_49_bF_buf0_), .Y(_17324_) );
OAI21X1 OAI21X1_2778 ( .gnd(gnd), .vdd(vdd), .A(_17323_), .B(_17324_), .C(_17273_), .Y(module_3_W_193_) );
AND2X2 AND2X2_404 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf4_), .B(bloque_datos_50_bF_buf1_), .Y(_17325_) );
NOR2X1 NOR2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf3_), .B(bloque_datos_50_bF_buf0_), .Y(_17326_) );
OAI21X1 OAI21X1_2779 ( .gnd(gnd), .vdd(vdd), .A(_17325_), .B(_17326_), .C(_17275_), .Y(module_3_W_194_) );
OR2X2 OR2X2_417 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_171_), .B(bloque_datos_51_bF_buf1_), .Y(module_3_W_195_) );
NOR2X1 NOR2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf1_), .B(module_3_W_172_), .Y(_17327_) );
INVX1 INVX1_2503 ( .gnd(gnd), .vdd(vdd), .A(_17327_), .Y(module_3_W_196_) );
NOR2X1 NOR2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf0_), .B(module_3_W_173_), .Y(_17328_) );
INVX1 INVX1_2504 ( .gnd(gnd), .vdd(vdd), .A(_17328_), .Y(module_3_W_197_) );
OR2X2 OR2X2_418 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_174_), .B(bloque_datos_54_bF_buf0_), .Y(module_3_W_198_) );
XNOR2X1 XNOR2X1_473 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf0_), .B(bloque_datos[55]), .Y(_17329_) );
NAND2X1 NAND2X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_17329_), .B(_17288_), .Y(module_3_W_199_) );
NAND2X1 NAND2X1_2303 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf2_), .B(module_3_W_128_), .Y(_17330_) );
INVX1 INVX1_2505 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf1_), .Y(_17331_) );
NAND2X1 NAND2X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_17331_), .B(_17228_), .Y(_17332_) );
AOI21X1 AOI21X1_2468 ( .gnd(gnd), .vdd(vdd), .A(_17332_), .B(_17330_), .C(module_3_W_176_), .Y(_17333_) );
INVX2 INVX2_618 ( .gnd(gnd), .vdd(vdd), .A(_17333_), .Y(module_3_W_200_) );
NAND2X1 NAND2X1_2305 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf1_), .B(module_3_W_129_), .Y(_17334_) );
OR2X2 OR2X2_419 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_129_), .B(bloque_datos_57_bF_buf0_), .Y(_17335_) );
AOI21X1 AOI21X1_2469 ( .gnd(gnd), .vdd(vdd), .A(_17334_), .B(_17335_), .C(module_3_W_177_), .Y(_17336_) );
INVX1 INVX1_2506 ( .gnd(gnd), .vdd(vdd), .A(_17336_), .Y(module_3_W_201_) );
NAND2X1 NAND2X1_2306 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf2_), .B(module_3_W_130_), .Y(_17337_) );
INVX1 INVX1_2507 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf1_), .Y(_17338_) );
NAND2X1 NAND2X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_17338_), .B(_17232_), .Y(_17339_) );
AOI21X1 AOI21X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_17339_), .B(_17337_), .C(module_3_W_178_), .Y(_17340_) );
INVX1 INVX1_2508 ( .gnd(gnd), .vdd(vdd), .A(_17340_), .Y(module_3_W_202_) );
NAND2X1 NAND2X1_2308 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf2_), .B(module_3_W_131_), .Y(_17341_) );
INVX1 INVX1_2509 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf1_), .Y(_17342_) );
NAND2X1 NAND2X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_17342_), .B(_17234_), .Y(_17343_) );
AOI21X1 AOI21X1_2471 ( .gnd(gnd), .vdd(vdd), .A(_17343_), .B(_17341_), .C(module_3_W_179_), .Y(_17344_) );
INVX1 INVX1_2510 ( .gnd(gnd), .vdd(vdd), .A(_17344_), .Y(module_3_W_203_) );
XNOR2X1 XNOR2X1_474 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_132_), .B(bloque_datos_60_bF_buf0_), .Y(_17345_) );
NAND2X1 NAND2X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_17345_), .B(_17298_), .Y(module_3_W_204_) );
NAND2X1 NAND2X1_2311 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf2_), .B(module_3_W_133_), .Y(_17346_) );
OR2X2 OR2X2_420 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_133_), .B(bloque_datos_61_bF_buf1_), .Y(_17347_) );
AOI21X1 AOI21X1_2472 ( .gnd(gnd), .vdd(vdd), .A(_17346_), .B(_17347_), .C(module_3_W_181_), .Y(_17348_) );
INVX1 INVX1_2511 ( .gnd(gnd), .vdd(vdd), .A(_17348_), .Y(module_3_W_205_) );
INVX2 INVX2_619 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf0_), .Y(_17349_) );
NAND2X1 NAND2X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_17349_), .B(_17306_), .Y(module_3_W_206_) );
INVX2 INVX2_620 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[63]), .Y(_17350_) );
NAND2X1 NAND2X1_2313 ( .gnd(gnd), .vdd(vdd), .A(_17350_), .B(_17308_), .Y(module_3_W_207_) );
OAI21X1 OAI21X1_2780 ( .gnd(gnd), .vdd(vdd), .A(_17248_), .B(bloque_datos_80_bF_buf5_), .C(bloque_datos_64_bF_buf2_), .Y(_17351_) );
OR2X2 OR2X2_421 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_136_), .B(bloque_datos_64_bF_buf1_), .Y(_17352_) );
AOI21X1 AOI21X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_17351_), .B(_17352_), .C(module_3_W_184_), .Y(_17353_) );
INVX1 INVX1_2512 ( .gnd(gnd), .vdd(vdd), .A(_17353_), .Y(module_3_W_208_) );
NAND2X1 NAND2X1_2314 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_65_bF_buf1_), .B(module_3_W_137_), .Y(_17354_) );
OR2X2 OR2X2_422 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_137_), .B(bloque_datos_65_bF_buf0_), .Y(_17355_) );
AOI21X1 AOI21X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_17354_), .B(_17355_), .C(module_3_W_185_), .Y(_17356_) );
INVX1 INVX1_2513 ( .gnd(gnd), .vdd(vdd), .A(_17356_), .Y(module_3_W_209_) );
OAI21X1 OAI21X1_2781 ( .gnd(gnd), .vdd(vdd), .A(_17256_), .B(bloque_datos_82_bF_buf3_), .C(bloque_datos_66_bF_buf2_), .Y(_17357_) );
OR2X2 OR2X2_423 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_138_), .B(bloque_datos_66_bF_buf1_), .Y(_17358_) );
AOI21X1 AOI21X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_17357_), .B(_17358_), .C(module_3_W_186_), .Y(_17359_) );
INVX1 INVX1_2514 ( .gnd(gnd), .vdd(vdd), .A(_17359_), .Y(module_3_W_210_) );
OAI21X1 OAI21X1_2782 ( .gnd(gnd), .vdd(vdd), .A(_17259_), .B(bloque_datos_83_bF_buf5_), .C(bloque_datos_67_bF_buf3_), .Y(_17360_) );
OR2X2 OR2X2_424 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_139_), .B(bloque_datos_67_bF_buf2_), .Y(_17361_) );
AOI21X1 AOI21X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_17360_), .B(_17361_), .C(module_3_W_187_), .Y(_17362_) );
INVX1 INVX1_2515 ( .gnd(gnd), .vdd(vdd), .A(_17362_), .Y(module_3_W_211_) );
NAND2X1 NAND2X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_17278_), .B(_17314_), .Y(module_3_W_212_) );
NAND2X1 NAND2X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_17281_), .B(_17316_), .Y(module_3_W_213_) );
NAND2X1 NAND2X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_17284_), .B(_17318_), .Y(module_3_W_214_) );
INVX1 INVX1_2516 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf0_), .Y(_17363_) );
NAND2X1 NAND2X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_17363_), .B(_17320_), .Y(module_3_W_215_) );
OR2X2 OR2X2_425 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_192_), .B(bloque_datos_72_bF_buf1_), .Y(module_3_W_216_) );
OR2X2 OR2X2_426 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_193_), .B(bloque_datos_73_bF_buf0_), .Y(module_3_W_217_) );
OR2X2 OR2X2_427 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_194_), .B(bloque_datos_74_bF_buf1_), .Y(module_3_W_218_) );
OR2X2 OR2X2_428 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_195_), .B(bloque_datos_75_bF_buf2_), .Y(module_3_W_219_) );
NAND2X1 NAND2X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_17237_), .B(_17327_), .Y(module_3_W_220_) );
NAND2X1 NAND2X1_2320 ( .gnd(gnd), .vdd(vdd), .A(_17300_), .B(_17328_), .Y(module_3_W_221_) );
OR2X2 OR2X2_429 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_198_), .B(bloque_datos_78_bF_buf1_), .Y(module_3_W_222_) );
OR2X2 OR2X2_430 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_199_), .B(bloque_datos_79_bF_buf0_), .Y(module_3_W_223_) );
XNOR2X1 XNOR2X1_475 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_152_), .B(bloque_datos_80_bF_buf4_), .Y(_17364_) );
NAND2X1 NAND2X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_17333_), .B(_17364_), .Y(module_3_W_224_) );
OAI21X1 OAI21X1_2783 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_129_), .B(_17230_), .C(bloque_datos_81_bF_buf1_), .Y(_17365_) );
NAND3X1 NAND3X1_3924 ( .gnd(gnd), .vdd(vdd), .A(_17252_), .B(_17293_), .C(_17292_), .Y(_17366_) );
NAND2X1 NAND2X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_17365_), .B(_17366_), .Y(_17367_) );
NAND2X1 NAND2X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_17367_), .B(_17336_), .Y(module_3_W_225_) );
XNOR2X1 XNOR2X1_476 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_154_), .B(bloque_datos_82_bF_buf2_), .Y(_17368_) );
NAND2X1 NAND2X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_17340_), .B(_17368_), .Y(module_3_W_226_) );
XNOR2X1 XNOR2X1_477 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_155_), .B(bloque_datos_83_bF_buf4_), .Y(_17369_) );
NAND2X1 NAND2X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_17344_), .B(_17369_), .Y(module_3_W_227_) );
INVX1 INVX1_2517 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf1_), .Y(_17370_) );
NAND3X1 NAND3X1_3925 ( .gnd(gnd), .vdd(vdd), .A(_17370_), .B(_17345_), .C(_17298_), .Y(module_3_W_228_) );
OAI21X1 OAI21X1_2784 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_133_), .B(_17242_), .C(bloque_datos_85_bF_buf3_), .Y(_17371_) );
INVX1 INVX1_2518 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf2_), .Y(_17372_) );
NAND3X1 NAND3X1_3926 ( .gnd(gnd), .vdd(vdd), .A(_17372_), .B(_17303_), .C(_17302_), .Y(_17373_) );
NAND2X1 NAND2X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_17371_), .B(_17373_), .Y(_17374_) );
NAND2X1 NAND2X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_17374_), .B(_17348_), .Y(module_3_W_229_) );
INVX1 INVX1_2519 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf1_), .Y(_17375_) );
NAND3X1 NAND3X1_3927 ( .gnd(gnd), .vdd(vdd), .A(_17375_), .B(_17349_), .C(_17306_), .Y(module_3_W_230_) );
INVX1 INVX1_2520 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf0_), .Y(_17376_) );
NAND3X1 NAND3X1_3928 ( .gnd(gnd), .vdd(vdd), .A(_17376_), .B(_17350_), .C(_17308_), .Y(module_3_W_231_) );
AOI21X1 AOI21X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_17250_), .B(_17249_), .C(_17197_), .Y(_17377_) );
NOR2X1 NOR2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf2_), .B(module_3_W_160_), .Y(_17378_) );
OAI21X1 OAI21X1_2785 ( .gnd(gnd), .vdd(vdd), .A(_17378_), .B(_17377_), .C(_17353_), .Y(module_3_W_232_) );
AOI21X1 AOI21X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_17255_), .B(_17254_), .C(_17201_), .Y(_17379_) );
NOR2X1 NOR2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf0_), .B(module_3_W_161_), .Y(_17380_) );
OAI21X1 OAI21X1_2786 ( .gnd(gnd), .vdd(vdd), .A(_17379_), .B(_17380_), .C(_17356_), .Y(module_3_W_233_) );
AOI21X1 AOI21X1_2479 ( .gnd(gnd), .vdd(vdd), .A(_17258_), .B(_17257_), .C(_17205_), .Y(_17381_) );
NOR2X1 NOR2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf2_), .B(module_3_W_162_), .Y(_17382_) );
OAI21X1 OAI21X1_2787 ( .gnd(gnd), .vdd(vdd), .A(_17382_), .B(_17381_), .C(_17359_), .Y(module_3_W_234_) );
AOI21X1 AOI21X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_17261_), .B(_17260_), .C(_17209_), .Y(_17383_) );
NOR2X1 NOR2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf0_), .B(module_3_W_163_), .Y(_17384_) );
OAI21X1 OAI21X1_2788 ( .gnd(gnd), .vdd(vdd), .A(_17384_), .B(_17383_), .C(_17362_), .Y(module_3_W_235_) );
NAND3X1 NAND3X1_3929 ( .gnd(gnd), .vdd(vdd), .A(_17213_), .B(_17278_), .C(_17314_), .Y(module_3_W_236_) );
NAND3X1 NAND3X1_3930 ( .gnd(gnd), .vdd(vdd), .A(_17217_), .B(_17281_), .C(_17316_), .Y(module_3_W_237_) );
NAND3X1 NAND3X1_3931 ( .gnd(gnd), .vdd(vdd), .A(_17221_), .B(_17284_), .C(_17318_), .Y(module_3_W_238_) );
NAND3X1 NAND3X1_3932 ( .gnd(gnd), .vdd(vdd), .A(_17225_), .B(_17363_), .C(_17320_), .Y(module_3_W_239_) );
OR2X2 OR2X2_431 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_192_), .B(module_3_W_128_), .Y(module_3_W_240_) );
OR2X2 OR2X2_432 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_193_), .B(module_3_W_129_), .Y(module_3_W_241_) );
OR2X2 OR2X2_433 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_194_), .B(module_3_W_130_), .Y(module_3_W_242_) );
OR2X2 OR2X2_434 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_195_), .B(module_3_W_131_), .Y(module_3_W_243_) );
NAND2X1 NAND2X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_17239_), .B(_17327_), .Y(module_3_W_244_) );
NAND2X1 NAND2X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_17302_), .B(_17328_), .Y(module_3_W_245_) );
OR2X2 OR2X2_435 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_198_), .B(module_3_W_134_), .Y(module_3_W_246_) );
OR2X2 OR2X2_436 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_199_), .B(module_3_W_135_), .Y(module_3_W_247_) );
XNOR2X1 XNOR2X1_478 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_176_), .B(module_3_W_136_), .Y(_17385_) );
NAND3X1 NAND3X1_3933 ( .gnd(gnd), .vdd(vdd), .A(_17333_), .B(_17364_), .C(_17385_), .Y(module_3_W_248_) );
NAND3X1 NAND3X1_3934 ( .gnd(gnd), .vdd(vdd), .A(_17254_), .B(_17367_), .C(_17336_), .Y(module_3_W_249_) );
XNOR2X1 XNOR2X1_479 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_178_), .B(module_3_W_138_), .Y(_17386_) );
NAND3X1 NAND3X1_3935 ( .gnd(gnd), .vdd(vdd), .A(_17340_), .B(_17368_), .C(_17386_), .Y(module_3_W_250_) );
XNOR2X1 XNOR2X1_480 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_179_), .B(module_3_W_139_), .Y(_17387_) );
NAND3X1 NAND3X1_3936 ( .gnd(gnd), .vdd(vdd), .A(_17344_), .B(_17369_), .C(_17387_), .Y(module_3_W_251_) );
INVX1 INVX1_2521 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_140_), .Y(_17388_) );
NAND3X1 NAND3X1_3937 ( .gnd(gnd), .vdd(vdd), .A(_17388_), .B(_17345_), .C(_17298_), .Y(module_3_W_252_) );
INVX1 INVX1_2522 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_141_), .Y(_17389_) );
NAND3X1 NAND3X1_3938 ( .gnd(gnd), .vdd(vdd), .A(_17389_), .B(_17374_), .C(_17348_), .Y(module_3_W_253_) );
INVX1 INVX1_2523 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_142_), .Y(_17390_) );
NAND3X1 NAND3X1_3939 ( .gnd(gnd), .vdd(vdd), .A(_17349_), .B(_17390_), .C(_17306_), .Y(module_3_W_254_) );
INVX1 INVX1_2524 ( .gnd(gnd), .vdd(vdd), .A(module_3_W_143_), .Y(_17391_) );
NAND3X1 NAND3X1_3940 ( .gnd(gnd), .vdd(vdd), .A(_17350_), .B(_17391_), .C(_17308_), .Y(module_3_W_255_) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(module_0_H_8_) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(module_0_H_9_) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(module_0_H_10_) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(module_0_H_11_) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(module_0_W_32_) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(module_0_W_33_) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf3_), .Y(module_0_W_34_) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf3_), .Y(module_0_W_35_) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf3_), .Y(module_0_W_36_) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf3_), .Y(module_0_W_37_) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf3_), .Y(module_0_W_38_) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[7]), .Y(module_0_W_39_) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .Y(module_0_W_40_) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .Y(module_0_W_41_) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .Y(module_0_W_42_) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .Y(module_0_W_43_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf3_), .Y(module_0_W_44_) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf3_), .Y(module_0_W_45_) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf3_), .Y(module_0_W_46_) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[15]), .Y(module_0_W_47_) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf3_), .Y(module_0_W_48_) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .Y(module_0_W_49_) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .Y(module_0_W_50_) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf3_), .Y(module_0_W_51_) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf3_), .Y(module_0_W_52_) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf3_), .Y(module_0_W_53_) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf3_), .Y(module_0_W_54_) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf3_), .Y(module_0_W_55_) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf0_), .Y(module_0_W_56_) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf3_), .Y(module_0_W_57_) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf3_), .Y(module_0_W_58_) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf1_), .Y(module_0_W_59_) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf1_), .Y(module_0_W_60_) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf1_), .Y(module_0_W_61_) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf3_), .Y(module_0_W_62_) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf3_), .Y(module_0_W_63_) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf0_), .Y(module_0_W_64_) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf3_), .Y(module_0_W_65_) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf0_), .Y(module_0_W_66_) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf0_), .Y(module_0_W_67_) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf3_), .Y(module_0_W_68_) );
BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf3_), .Y(module_0_W_69_) );
BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf3_), .Y(module_0_W_70_) );
BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .Y(module_0_W_71_) );
BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf0_), .Y(module_0_W_72_) );
BUFX2 BUFX2_71 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf3_), .Y(module_0_W_73_) );
BUFX2 BUFX2_72 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf3_), .Y(module_0_W_74_) );
BUFX2 BUFX2_73 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf3_), .Y(module_0_W_75_) );
BUFX2 BUFX2_74 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf0_), .Y(module_0_W_76_) );
BUFX2 BUFX2_75 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf0_), .Y(module_0_W_77_) );
BUFX2 BUFX2_76 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf0_), .Y(module_0_W_78_) );
BUFX2 BUFX2_77 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_47_bF_buf3_), .Y(module_0_W_79_) );
BUFX2 BUFX2_78 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_48_bF_buf0_), .Y(module_0_W_80_) );
BUFX2 BUFX2_79 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_49_bF_buf3_), .Y(module_0_W_81_) );
BUFX2 BUFX2_80 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_50_bF_buf3_), .Y(module_0_W_82_) );
BUFX2 BUFX2_81 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf0_), .Y(module_0_W_83_) );
BUFX2 BUFX2_82 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf0_), .Y(module_0_W_84_) );
BUFX2 BUFX2_83 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf3_), .Y(module_0_W_85_) );
BUFX2 BUFX2_84 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf3_), .Y(module_0_W_86_) );
BUFX2 BUFX2_85 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[55]), .Y(module_0_W_87_) );
BUFX2 BUFX2_86 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf0_), .Y(module_0_W_88_) );
BUFX2 BUFX2_87 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf3_), .Y(module_0_W_89_) );
BUFX2 BUFX2_88 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf0_), .Y(module_0_W_90_) );
BUFX2 BUFX2_89 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf0_), .Y(module_0_W_91_) );
BUFX2 BUFX2_90 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf3_), .Y(module_0_W_92_) );
BUFX2 BUFX2_91 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf0_), .Y(module_0_W_93_) );
BUFX2 BUFX2_92 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf3_), .Y(module_0_W_94_) );
BUFX2 BUFX2_93 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[63]), .Y(module_0_W_95_) );
BUFX2 BUFX2_94 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_64_bF_buf0_), .Y(module_0_W_96_) );
BUFX2 BUFX2_95 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_65_bF_buf3_), .Y(module_0_W_97_) );
BUFX2 BUFX2_96 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf0_), .Y(module_0_W_98_) );
BUFX2 BUFX2_97 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf1_), .Y(module_0_W_99_) );
BUFX2 BUFX2_98 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf3_), .Y(module_0_W_100_) );
BUFX2 BUFX2_99 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf3_), .Y(module_0_W_101_) );
BUFX2 BUFX2_100 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf3_), .Y(module_0_W_102_) );
BUFX2 BUFX2_101 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf3_), .Y(module_0_W_103_) );
BUFX2 BUFX2_102 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf0_), .Y(module_0_W_104_) );
BUFX2 BUFX2_103 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_73_bF_buf3_), .Y(module_0_W_105_) );
BUFX2 BUFX2_104 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf0_), .Y(module_0_W_106_) );
BUFX2 BUFX2_105 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf1_), .Y(module_0_W_107_) );
BUFX2 BUFX2_106 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf0_), .Y(module_0_W_108_) );
BUFX2 BUFX2_107 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf0_), .Y(module_0_W_109_) );
BUFX2 BUFX2_108 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf0_), .Y(module_0_W_110_) );
BUFX2 BUFX2_109 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_79_bF_buf3_), .Y(module_0_W_111_) );
BUFX2 BUFX2_110 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf3_), .Y(module_0_W_112_) );
BUFX2 BUFX2_111 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf0_), .Y(module_0_W_113_) );
BUFX2 BUFX2_112 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf1_), .Y(module_0_W_114_) );
BUFX2 BUFX2_113 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf3_), .Y(module_0_W_115_) );
BUFX2 BUFX2_114 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf0_), .Y(module_0_W_116_) );
BUFX2 BUFX2_115 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf1_), .Y(module_0_W_117_) );
BUFX2 BUFX2_116 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf0_), .Y(module_0_W_118_) );
BUFX2 BUFX2_117 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf3_), .Y(module_0_W_119_) );
BUFX2 BUFX2_118 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf1_), .Y(module_0_W_120_) );
BUFX2 BUFX2_119 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf3_), .Y(module_0_W_121_) );
BUFX2 BUFX2_120 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf1_), .Y(module_0_W_122_) );
BUFX2 BUFX2_121 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf3_), .Y(module_0_W_123_) );
BUFX2 BUFX2_122 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf3_), .Y(module_0_W_124_) );
BUFX2 BUFX2_123 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf3_), .Y(module_0_W_125_) );
BUFX2 BUFX2_124 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf3_), .Y(module_0_W_126_) );
BUFX2 BUFX2_125 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf3_), .Y(module_0_W_127_) );
BUFX2 BUFX2_126 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(module_1_H_8_) );
BUFX2 BUFX2_127 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(module_1_H_9_) );
BUFX2 BUFX2_128 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(module_1_H_10_) );
BUFX2 BUFX2_129 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(module_1_H_11_) );
BUFX2 BUFX2_130 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(module_1_W_32_) );
BUFX2 BUFX2_131 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(module_1_W_33_) );
BUFX2 BUFX2_132 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf2_), .Y(module_1_W_34_) );
BUFX2 BUFX2_133 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf2_), .Y(module_1_W_35_) );
BUFX2 BUFX2_134 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf2_), .Y(module_1_W_36_) );
BUFX2 BUFX2_135 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf2_), .Y(module_1_W_37_) );
BUFX2 BUFX2_136 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf2_), .Y(module_1_W_38_) );
BUFX2 BUFX2_137 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[7]), .Y(module_1_W_39_) );
BUFX2 BUFX2_138 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .Y(module_1_W_40_) );
BUFX2 BUFX2_139 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .Y(module_1_W_41_) );
BUFX2 BUFX2_140 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .Y(module_1_W_42_) );
BUFX2 BUFX2_141 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .Y(module_1_W_43_) );
BUFX2 BUFX2_142 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf2_), .Y(module_1_W_44_) );
BUFX2 BUFX2_143 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf2_), .Y(module_1_W_45_) );
BUFX2 BUFX2_144 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf2_), .Y(module_1_W_46_) );
BUFX2 BUFX2_145 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[15]), .Y(module_1_W_47_) );
BUFX2 BUFX2_146 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf2_), .Y(module_1_W_48_) );
BUFX2 BUFX2_147 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .Y(module_1_W_49_) );
BUFX2 BUFX2_148 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .Y(module_1_W_50_) );
BUFX2 BUFX2_149 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf2_), .Y(module_1_W_51_) );
BUFX2 BUFX2_150 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf2_), .Y(module_1_W_52_) );
BUFX2 BUFX2_151 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf2_), .Y(module_1_W_53_) );
BUFX2 BUFX2_152 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf2_), .Y(module_1_W_54_) );
BUFX2 BUFX2_153 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf2_), .Y(module_1_W_55_) );
BUFX2 BUFX2_154 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf4_), .Y(module_1_W_56_) );
BUFX2 BUFX2_155 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf2_), .Y(module_1_W_57_) );
BUFX2 BUFX2_156 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf2_), .Y(module_1_W_58_) );
BUFX2 BUFX2_157 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf0_), .Y(module_1_W_59_) );
BUFX2 BUFX2_158 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf0_), .Y(module_1_W_60_) );
BUFX2 BUFX2_159 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf0_), .Y(module_1_W_61_) );
BUFX2 BUFX2_160 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf2_), .Y(module_1_W_62_) );
BUFX2 BUFX2_161 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf2_), .Y(module_1_W_63_) );
BUFX2 BUFX2_162 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf4_), .Y(module_1_W_64_) );
BUFX2 BUFX2_163 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf2_), .Y(module_1_W_65_) );
BUFX2 BUFX2_164 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf4_), .Y(module_1_W_66_) );
BUFX2 BUFX2_165 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf4_), .Y(module_1_W_67_) );
BUFX2 BUFX2_166 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf2_), .Y(module_1_W_68_) );
BUFX2 BUFX2_167 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf2_), .Y(module_1_W_69_) );
BUFX2 BUFX2_168 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf2_), .Y(module_1_W_70_) );
BUFX2 BUFX2_169 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .Y(module_1_W_71_) );
BUFX2 BUFX2_170 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf4_), .Y(module_1_W_72_) );
BUFX2 BUFX2_171 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf2_), .Y(module_1_W_73_) );
BUFX2 BUFX2_172 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf2_), .Y(module_1_W_74_) );
BUFX2 BUFX2_173 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf2_), .Y(module_1_W_75_) );
BUFX2 BUFX2_174 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf4_), .Y(module_1_W_76_) );
BUFX2 BUFX2_175 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf4_), .Y(module_1_W_77_) );
BUFX2 BUFX2_176 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf4_), .Y(module_1_W_78_) );
BUFX2 BUFX2_177 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_47_bF_buf2_), .Y(module_1_W_79_) );
BUFX2 BUFX2_178 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_48_bF_buf4_), .Y(module_1_W_80_) );
BUFX2 BUFX2_179 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_49_bF_buf2_), .Y(module_1_W_81_) );
BUFX2 BUFX2_180 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_50_bF_buf2_), .Y(module_1_W_82_) );
BUFX2 BUFX2_181 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf4_), .Y(module_1_W_83_) );
BUFX2 BUFX2_182 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf4_), .Y(module_1_W_84_) );
BUFX2 BUFX2_183 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf2_), .Y(module_1_W_85_) );
BUFX2 BUFX2_184 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf2_), .Y(module_1_W_86_) );
BUFX2 BUFX2_185 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[55]), .Y(module_1_W_87_) );
BUFX2 BUFX2_186 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf4_), .Y(module_1_W_88_) );
BUFX2 BUFX2_187 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf2_), .Y(module_1_W_89_) );
BUFX2 BUFX2_188 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf4_), .Y(module_1_W_90_) );
BUFX2 BUFX2_189 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf4_), .Y(module_1_W_91_) );
BUFX2 BUFX2_190 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf2_), .Y(module_1_W_92_) );
BUFX2 BUFX2_191 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf4_), .Y(module_1_W_93_) );
BUFX2 BUFX2_192 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf2_), .Y(module_1_W_94_) );
BUFX2 BUFX2_193 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[63]), .Y(module_1_W_95_) );
BUFX2 BUFX2_194 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_64_bF_buf4_), .Y(module_1_W_96_) );
BUFX2 BUFX2_195 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_65_bF_buf2_), .Y(module_1_W_97_) );
BUFX2 BUFX2_196 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf4_), .Y(module_1_W_98_) );
BUFX2 BUFX2_197 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf0_), .Y(module_1_W_99_) );
BUFX2 BUFX2_198 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf2_), .Y(module_1_W_100_) );
BUFX2 BUFX2_199 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf2_), .Y(module_1_W_101_) );
BUFX2 BUFX2_200 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf2_), .Y(module_1_W_102_) );
BUFX2 BUFX2_201 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf2_), .Y(module_1_W_103_) );
BUFX2 BUFX2_202 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf4_), .Y(module_1_W_104_) );
BUFX2 BUFX2_203 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_73_bF_buf2_), .Y(module_1_W_105_) );
BUFX2 BUFX2_204 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf4_), .Y(module_1_W_106_) );
BUFX2 BUFX2_205 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf0_), .Y(module_1_W_107_) );
BUFX2 BUFX2_206 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf4_), .Y(module_1_W_108_) );
BUFX2 BUFX2_207 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf4_), .Y(module_1_W_109_) );
BUFX2 BUFX2_208 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf4_), .Y(module_1_W_110_) );
BUFX2 BUFX2_209 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_79_bF_buf2_), .Y(module_1_W_111_) );
BUFX2 BUFX2_210 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf2_), .Y(module_1_W_112_) );
BUFX2 BUFX2_211 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf4_), .Y(module_1_W_113_) );
BUFX2 BUFX2_212 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf0_), .Y(module_1_W_114_) );
BUFX2 BUFX2_213 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf2_), .Y(module_1_W_115_) );
BUFX2 BUFX2_214 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf4_), .Y(module_1_W_116_) );
BUFX2 BUFX2_215 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf0_), .Y(module_1_W_117_) );
BUFX2 BUFX2_216 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf4_), .Y(module_1_W_118_) );
BUFX2 BUFX2_217 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf2_), .Y(module_1_W_119_) );
BUFX2 BUFX2_218 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf0_), .Y(module_1_W_120_) );
BUFX2 BUFX2_219 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf2_), .Y(module_1_W_121_) );
BUFX2 BUFX2_220 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf0_), .Y(module_1_W_122_) );
BUFX2 BUFX2_221 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf2_), .Y(module_1_W_123_) );
BUFX2 BUFX2_222 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf2_), .Y(module_1_W_124_) );
BUFX2 BUFX2_223 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf2_), .Y(module_1_W_125_) );
BUFX2 BUFX2_224 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf2_), .Y(module_1_W_126_) );
BUFX2 BUFX2_225 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf2_), .Y(module_1_W_127_) );
BUFX2 BUFX2_226 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(module_2_H_8_) );
BUFX2 BUFX2_227 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(module_2_H_9_) );
BUFX2 BUFX2_228 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(module_2_H_10_) );
BUFX2 BUFX2_229 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(module_2_H_11_) );
BUFX2 BUFX2_230 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(module_2_W_32_) );
BUFX2 BUFX2_231 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(module_2_W_33_) );
BUFX2 BUFX2_232 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf1_), .Y(module_2_W_34_) );
BUFX2 BUFX2_233 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf1_), .Y(module_2_W_35_) );
BUFX2 BUFX2_234 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf1_), .Y(module_2_W_36_) );
BUFX2 BUFX2_235 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf1_), .Y(module_2_W_37_) );
BUFX2 BUFX2_236 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf1_), .Y(module_2_W_38_) );
BUFX2 BUFX2_237 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[7]), .Y(module_2_W_39_) );
BUFX2 BUFX2_238 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .Y(module_2_W_40_) );
BUFX2 BUFX2_239 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .Y(module_2_W_41_) );
BUFX2 BUFX2_240 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .Y(module_2_W_42_) );
BUFX2 BUFX2_241 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .Y(module_2_W_43_) );
BUFX2 BUFX2_242 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf1_), .Y(module_2_W_44_) );
BUFX2 BUFX2_243 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf1_), .Y(module_2_W_45_) );
BUFX2 BUFX2_244 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf1_), .Y(module_2_W_46_) );
BUFX2 BUFX2_245 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[15]), .Y(module_2_W_47_) );
BUFX2 BUFX2_246 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf1_), .Y(module_2_W_48_) );
BUFX2 BUFX2_247 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .Y(module_2_W_49_) );
BUFX2 BUFX2_248 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .Y(module_2_W_50_) );
BUFX2 BUFX2_249 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf1_), .Y(module_2_W_51_) );
BUFX2 BUFX2_250 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf1_), .Y(module_2_W_52_) );
BUFX2 BUFX2_251 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf1_), .Y(module_2_W_53_) );
BUFX2 BUFX2_252 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf1_), .Y(module_2_W_54_) );
BUFX2 BUFX2_253 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf1_), .Y(module_2_W_55_) );
BUFX2 BUFX2_254 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf3_), .Y(module_2_W_56_) );
BUFX2 BUFX2_255 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf1_), .Y(module_2_W_57_) );
BUFX2 BUFX2_256 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf1_), .Y(module_2_W_58_) );
BUFX2 BUFX2_257 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf4_), .Y(module_2_W_59_) );
BUFX2 BUFX2_258 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf4_), .Y(module_2_W_60_) );
BUFX2 BUFX2_259 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf4_), .Y(module_2_W_61_) );
BUFX2 BUFX2_260 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf1_), .Y(module_2_W_62_) );
BUFX2 BUFX2_261 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf1_), .Y(module_2_W_63_) );
BUFX2 BUFX2_262 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf3_), .Y(module_2_W_64_) );
BUFX2 BUFX2_263 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf1_), .Y(module_2_W_65_) );
BUFX2 BUFX2_264 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf3_), .Y(module_2_W_66_) );
BUFX2 BUFX2_265 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf3_), .Y(module_2_W_67_) );
BUFX2 BUFX2_266 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf1_), .Y(module_2_W_68_) );
BUFX2 BUFX2_267 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf1_), .Y(module_2_W_69_) );
BUFX2 BUFX2_268 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf1_), .Y(module_2_W_70_) );
BUFX2 BUFX2_269 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .Y(module_2_W_71_) );
BUFX2 BUFX2_270 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf3_), .Y(module_2_W_72_) );
BUFX2 BUFX2_271 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf1_), .Y(module_2_W_73_) );
BUFX2 BUFX2_272 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf1_), .Y(module_2_W_74_) );
BUFX2 BUFX2_273 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf1_), .Y(module_2_W_75_) );
BUFX2 BUFX2_274 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf3_), .Y(module_2_W_76_) );
BUFX2 BUFX2_275 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf3_), .Y(module_2_W_77_) );
BUFX2 BUFX2_276 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf3_), .Y(module_2_W_78_) );
BUFX2 BUFX2_277 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_47_bF_buf1_), .Y(module_2_W_79_) );
BUFX2 BUFX2_278 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_48_bF_buf3_), .Y(module_2_W_80_) );
BUFX2 BUFX2_279 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_49_bF_buf1_), .Y(module_2_W_81_) );
BUFX2 BUFX2_280 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_50_bF_buf1_), .Y(module_2_W_82_) );
BUFX2 BUFX2_281 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf3_), .Y(module_2_W_83_) );
BUFX2 BUFX2_282 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf3_), .Y(module_2_W_84_) );
BUFX2 BUFX2_283 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf1_), .Y(module_2_W_85_) );
BUFX2 BUFX2_284 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf1_), .Y(module_2_W_86_) );
BUFX2 BUFX2_285 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[55]), .Y(module_2_W_87_) );
BUFX2 BUFX2_286 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf3_), .Y(module_2_W_88_) );
BUFX2 BUFX2_287 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf1_), .Y(module_2_W_89_) );
BUFX2 BUFX2_288 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf3_), .Y(module_2_W_90_) );
BUFX2 BUFX2_289 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf3_), .Y(module_2_W_91_) );
BUFX2 BUFX2_290 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf1_), .Y(module_2_W_92_) );
BUFX2 BUFX2_291 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf3_), .Y(module_2_W_93_) );
BUFX2 BUFX2_292 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf1_), .Y(module_2_W_94_) );
BUFX2 BUFX2_293 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[63]), .Y(module_2_W_95_) );
BUFX2 BUFX2_294 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_64_bF_buf3_), .Y(module_2_W_96_) );
BUFX2 BUFX2_295 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_65_bF_buf1_), .Y(module_2_W_97_) );
BUFX2 BUFX2_296 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf3_), .Y(module_2_W_98_) );
BUFX2 BUFX2_297 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf4_), .Y(module_2_W_99_) );
BUFX2 BUFX2_298 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf1_), .Y(module_2_W_100_) );
BUFX2 BUFX2_299 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf1_), .Y(module_2_W_101_) );
BUFX2 BUFX2_300 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf1_), .Y(module_2_W_102_) );
BUFX2 BUFX2_301 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf1_), .Y(module_2_W_103_) );
BUFX2 BUFX2_302 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf3_), .Y(module_2_W_104_) );
BUFX2 BUFX2_303 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_73_bF_buf1_), .Y(module_2_W_105_) );
BUFX2 BUFX2_304 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf3_), .Y(module_2_W_106_) );
BUFX2 BUFX2_305 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf4_), .Y(module_2_W_107_) );
BUFX2 BUFX2_306 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf3_), .Y(module_2_W_108_) );
BUFX2 BUFX2_307 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf3_), .Y(module_2_W_109_) );
BUFX2 BUFX2_308 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf3_), .Y(module_2_W_110_) );
BUFX2 BUFX2_309 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_79_bF_buf1_), .Y(module_2_W_111_) );
BUFX2 BUFX2_310 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf1_), .Y(module_2_W_112_) );
BUFX2 BUFX2_311 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf3_), .Y(module_2_W_113_) );
BUFX2 BUFX2_312 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf4_), .Y(module_2_W_114_) );
BUFX2 BUFX2_313 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf1_), .Y(module_2_W_115_) );
BUFX2 BUFX2_314 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf3_), .Y(module_2_W_116_) );
BUFX2 BUFX2_315 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf4_), .Y(module_2_W_117_) );
BUFX2 BUFX2_316 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf3_), .Y(module_2_W_118_) );
BUFX2 BUFX2_317 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf1_), .Y(module_2_W_119_) );
BUFX2 BUFX2_318 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf4_), .Y(module_2_W_120_) );
BUFX2 BUFX2_319 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf1_), .Y(module_2_W_121_) );
BUFX2 BUFX2_320 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf4_), .Y(module_2_W_122_) );
BUFX2 BUFX2_321 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf1_), .Y(module_2_W_123_) );
BUFX2 BUFX2_322 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf1_), .Y(module_2_W_124_) );
BUFX2 BUFX2_323 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf1_), .Y(module_2_W_125_) );
BUFX2 BUFX2_324 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf1_), .Y(module_2_W_126_) );
BUFX2 BUFX2_325 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf1_), .Y(module_2_W_127_) );
BUFX2 BUFX2_326 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(module_3_H_8_) );
BUFX2 BUFX2_327 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(module_3_H_9_) );
BUFX2 BUFX2_328 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(module_3_H_10_) );
BUFX2 BUFX2_329 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(module_3_H_11_) );
BUFX2 BUFX2_330 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[0]), .Y(module_3_W_32_) );
BUFX2 BUFX2_331 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[1]), .Y(module_3_W_33_) );
BUFX2 BUFX2_332 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_2_bF_buf0_), .Y(module_3_W_34_) );
BUFX2 BUFX2_333 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_3_bF_buf0_), .Y(module_3_W_35_) );
BUFX2 BUFX2_334 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_4_bF_buf0_), .Y(module_3_W_36_) );
BUFX2 BUFX2_335 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_5_bF_buf0_), .Y(module_3_W_37_) );
BUFX2 BUFX2_336 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_6_bF_buf0_), .Y(module_3_W_38_) );
BUFX2 BUFX2_337 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[7]), .Y(module_3_W_39_) );
BUFX2 BUFX2_338 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[8]), .Y(module_3_W_40_) );
BUFX2 BUFX2_339 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[9]), .Y(module_3_W_41_) );
BUFX2 BUFX2_340 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[10]), .Y(module_3_W_42_) );
BUFX2 BUFX2_341 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[11]), .Y(module_3_W_43_) );
BUFX2 BUFX2_342 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_12_bF_buf0_), .Y(module_3_W_44_) );
BUFX2 BUFX2_343 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_13_bF_buf0_), .Y(module_3_W_45_) );
BUFX2 BUFX2_344 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_14_bF_buf0_), .Y(module_3_W_46_) );
BUFX2 BUFX2_345 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[15]), .Y(module_3_W_47_) );
BUFX2 BUFX2_346 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_16_bF_buf0_), .Y(module_3_W_48_) );
BUFX2 BUFX2_347 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[17]), .Y(module_3_W_49_) );
BUFX2 BUFX2_348 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[18]), .Y(module_3_W_50_) );
BUFX2 BUFX2_349 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_19_bF_buf0_), .Y(module_3_W_51_) );
BUFX2 BUFX2_350 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_20_bF_buf0_), .Y(module_3_W_52_) );
BUFX2 BUFX2_351 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_21_bF_buf0_), .Y(module_3_W_53_) );
BUFX2 BUFX2_352 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_22_bF_buf0_), .Y(module_3_W_54_) );
BUFX2 BUFX2_353 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_23_bF_buf0_), .Y(module_3_W_55_) );
BUFX2 BUFX2_354 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_24_bF_buf2_), .Y(module_3_W_56_) );
BUFX2 BUFX2_355 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_25_bF_buf0_), .Y(module_3_W_57_) );
BUFX2 BUFX2_356 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_26_bF_buf0_), .Y(module_3_W_58_) );
BUFX2 BUFX2_357 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_27_bF_buf3_), .Y(module_3_W_59_) );
BUFX2 BUFX2_358 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_28_bF_buf3_), .Y(module_3_W_60_) );
BUFX2 BUFX2_359 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_29_bF_buf3_), .Y(module_3_W_61_) );
BUFX2 BUFX2_360 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_30_bF_buf0_), .Y(module_3_W_62_) );
BUFX2 BUFX2_361 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_31_bF_buf0_), .Y(module_3_W_63_) );
BUFX2 BUFX2_362 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_32_bF_buf2_), .Y(module_3_W_64_) );
BUFX2 BUFX2_363 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_33_bF_buf0_), .Y(module_3_W_65_) );
BUFX2 BUFX2_364 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_34_bF_buf2_), .Y(module_3_W_66_) );
BUFX2 BUFX2_365 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_35_bF_buf2_), .Y(module_3_W_67_) );
BUFX2 BUFX2_366 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_36_bF_buf0_), .Y(module_3_W_68_) );
BUFX2 BUFX2_367 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_37_bF_buf0_), .Y(module_3_W_69_) );
BUFX2 BUFX2_368 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_38_bF_buf0_), .Y(module_3_W_70_) );
BUFX2 BUFX2_369 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[39]), .Y(module_3_W_71_) );
BUFX2 BUFX2_370 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_40_bF_buf2_), .Y(module_3_W_72_) );
BUFX2 BUFX2_371 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_41_bF_buf0_), .Y(module_3_W_73_) );
BUFX2 BUFX2_372 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_42_bF_buf0_), .Y(module_3_W_74_) );
BUFX2 BUFX2_373 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_43_bF_buf0_), .Y(module_3_W_75_) );
BUFX2 BUFX2_374 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_44_bF_buf2_), .Y(module_3_W_76_) );
BUFX2 BUFX2_375 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_45_bF_buf2_), .Y(module_3_W_77_) );
BUFX2 BUFX2_376 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_46_bF_buf2_), .Y(module_3_W_78_) );
BUFX2 BUFX2_377 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_47_bF_buf0_), .Y(module_3_W_79_) );
BUFX2 BUFX2_378 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_48_bF_buf2_), .Y(module_3_W_80_) );
BUFX2 BUFX2_379 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_49_bF_buf0_), .Y(module_3_W_81_) );
BUFX2 BUFX2_380 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_50_bF_buf0_), .Y(module_3_W_82_) );
BUFX2 BUFX2_381 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_51_bF_buf2_), .Y(module_3_W_83_) );
BUFX2 BUFX2_382 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_52_bF_buf2_), .Y(module_3_W_84_) );
BUFX2 BUFX2_383 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_53_bF_buf0_), .Y(module_3_W_85_) );
BUFX2 BUFX2_384 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_54_bF_buf0_), .Y(module_3_W_86_) );
BUFX2 BUFX2_385 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[55]), .Y(module_3_W_87_) );
BUFX2 BUFX2_386 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_56_bF_buf2_), .Y(module_3_W_88_) );
BUFX2 BUFX2_387 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_57_bF_buf0_), .Y(module_3_W_89_) );
BUFX2 BUFX2_388 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_58_bF_buf2_), .Y(module_3_W_90_) );
BUFX2 BUFX2_389 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_59_bF_buf2_), .Y(module_3_W_91_) );
BUFX2 BUFX2_390 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_60_bF_buf0_), .Y(module_3_W_92_) );
BUFX2 BUFX2_391 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_61_bF_buf2_), .Y(module_3_W_93_) );
BUFX2 BUFX2_392 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_62_bF_buf0_), .Y(module_3_W_94_) );
BUFX2 BUFX2_393 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos[63]), .Y(module_3_W_95_) );
BUFX2 BUFX2_394 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_64_bF_buf2_), .Y(module_3_W_96_) );
BUFX2 BUFX2_395 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_65_bF_buf0_), .Y(module_3_W_97_) );
BUFX2 BUFX2_396 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_66_bF_buf2_), .Y(module_3_W_98_) );
BUFX2 BUFX2_397 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_67_bF_buf3_), .Y(module_3_W_99_) );
BUFX2 BUFX2_398 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_68_bF_buf0_), .Y(module_3_W_100_) );
BUFX2 BUFX2_399 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_69_bF_buf0_), .Y(module_3_W_101_) );
BUFX2 BUFX2_400 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_70_bF_buf0_), .Y(module_3_W_102_) );
BUFX2 BUFX2_401 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_71_bF_buf0_), .Y(module_3_W_103_) );
BUFX2 BUFX2_402 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_72_bF_buf2_), .Y(module_3_W_104_) );
BUFX2 BUFX2_403 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_73_bF_buf0_), .Y(module_3_W_105_) );
BUFX2 BUFX2_404 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_74_bF_buf2_), .Y(module_3_W_106_) );
BUFX2 BUFX2_405 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_75_bF_buf3_), .Y(module_3_W_107_) );
BUFX2 BUFX2_406 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_76_bF_buf2_), .Y(module_3_W_108_) );
BUFX2 BUFX2_407 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_77_bF_buf2_), .Y(module_3_W_109_) );
BUFX2 BUFX2_408 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_78_bF_buf2_), .Y(module_3_W_110_) );
BUFX2 BUFX2_409 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_79_bF_buf0_), .Y(module_3_W_111_) );
BUFX2 BUFX2_410 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_80_bF_buf0_), .Y(module_3_W_112_) );
BUFX2 BUFX2_411 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_81_bF_buf2_), .Y(module_3_W_113_) );
BUFX2 BUFX2_412 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_82_bF_buf3_), .Y(module_3_W_114_) );
BUFX2 BUFX2_413 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_83_bF_buf0_), .Y(module_3_W_115_) );
BUFX2 BUFX2_414 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_84_bF_buf2_), .Y(module_3_W_116_) );
BUFX2 BUFX2_415 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_85_bF_buf3_), .Y(module_3_W_117_) );
BUFX2 BUFX2_416 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_86_bF_buf2_), .Y(module_3_W_118_) );
BUFX2 BUFX2_417 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_87_bF_buf0_), .Y(module_3_W_119_) );
BUFX2 BUFX2_418 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_88_bF_buf3_), .Y(module_3_W_120_) );
BUFX2 BUFX2_419 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_89_bF_buf0_), .Y(module_3_W_121_) );
BUFX2 BUFX2_420 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_90_bF_buf3_), .Y(module_3_W_122_) );
BUFX2 BUFX2_421 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_91_bF_buf0_), .Y(module_3_W_123_) );
BUFX2 BUFX2_422 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_92_bF_buf0_), .Y(module_3_W_124_) );
BUFX2 BUFX2_423 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_93_bF_buf0_), .Y(module_3_W_125_) );
BUFX2 BUFX2_424 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_94_bF_buf0_), .Y(module_3_W_126_) );
BUFX2 BUFX2_425 ( .gnd(gnd), .vdd(vdd), .A(bloque_datos_95_bF_buf0_), .Y(module_3_W_127_) );
endmodule
